
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"c1",x"c3",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"d8",x"c1",x"c3"),
    18 => (x"48",x"f4",x"e9",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"f4",x"e9",x"c2",x"87"),
    25 => (x"f0",x"e9",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"ef",x"c1",x"87",x"f7"),
    29 => (x"e9",x"c2",x"87",x"ee"),
    30 => (x"e9",x"c2",x"4d",x"f4"),
    31 => (x"ad",x"74",x"4c",x"f4"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"d0",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"c3",x"4c",x"87",x"ca"),
    69 => (x"74",x"9c",x"98",x"df"),
    70 => (x"87",x"eb",x"02",x"88"),
    71 => (x"4b",x"26",x"4a",x"26"),
    72 => (x"4f",x"26",x"4c",x"26"),
    73 => (x"81",x"48",x"73",x"1e"),
    74 => (x"c5",x"02",x"a9",x"73"),
    75 => (x"05",x"53",x"12",x"87"),
    76 => (x"4f",x"26",x"87",x"f6"),
    77 => (x"72",x"1e",x"73",x"1e"),
    78 => (x"e7",x"c0",x"02",x"9a"),
    79 => (x"c1",x"48",x"c0",x"87"),
    80 => (x"06",x"a9",x"72",x"4b"),
    81 => (x"82",x"72",x"87",x"d1"),
    82 => (x"73",x"87",x"c9",x"06"),
    83 => (x"01",x"a9",x"72",x"83"),
    84 => (x"87",x"c3",x"87",x"f4"),
    85 => (x"72",x"3a",x"b2",x"c1"),
    86 => (x"73",x"89",x"03",x"a9"),
    87 => (x"2a",x"c1",x"07",x"80"),
    88 => (x"87",x"f3",x"05",x"2b"),
    89 => (x"4f",x"26",x"4b",x"26"),
    90 => (x"c4",x"1e",x"75",x"1e"),
    91 => (x"a1",x"b7",x"71",x"4d"),
    92 => (x"c1",x"b9",x"ff",x"04"),
    93 => (x"07",x"bd",x"c3",x"81"),
    94 => (x"04",x"a2",x"b7",x"72"),
    95 => (x"82",x"c1",x"ba",x"ff"),
    96 => (x"fe",x"07",x"bd",x"c1"),
    97 => (x"2d",x"c1",x"87",x"ee"),
    98 => (x"c1",x"b8",x"ff",x"04"),
    99 => (x"04",x"2d",x"07",x"80"),
   100 => (x"81",x"c1",x"b9",x"ff"),
   101 => (x"26",x"4d",x"26",x"07"),
   102 => (x"1e",x"73",x"1e",x"4f"),
   103 => (x"66",x"c8",x"4a",x"71"),
   104 => (x"8b",x"c1",x"49",x"4b"),
   105 => (x"cf",x"02",x"99",x"71"),
   106 => (x"ff",x"48",x"12",x"87"),
   107 => (x"73",x"78",x"08",x"d4"),
   108 => (x"71",x"8b",x"c1",x"49"),
   109 => (x"87",x"f1",x"05",x"99"),
   110 => (x"4f",x"26",x"4b",x"26"),
   111 => (x"5c",x"5b",x"5e",x"0e"),
   112 => (x"ff",x"4a",x"71",x"0e"),
   113 => (x"66",x"cc",x"4c",x"d4"),
   114 => (x"8b",x"c1",x"49",x"4b"),
   115 => (x"ce",x"02",x"99",x"71"),
   116 => (x"7c",x"ff",x"c3",x"87"),
   117 => (x"49",x"73",x"52",x"6c"),
   118 => (x"99",x"71",x"8b",x"c1"),
   119 => (x"26",x"87",x"f2",x"05"),
   120 => (x"26",x"4b",x"26",x"4c"),
   121 => (x"1e",x"73",x"1e",x"4f"),
   122 => (x"c3",x"4b",x"d4",x"ff"),
   123 => (x"4a",x"6b",x"7b",x"ff"),
   124 => (x"6b",x"7b",x"ff",x"c3"),
   125 => (x"72",x"32",x"c8",x"49"),
   126 => (x"7b",x"ff",x"c3",x"b1"),
   127 => (x"31",x"c8",x"4a",x"6b"),
   128 => (x"ff",x"c3",x"b2",x"71"),
   129 => (x"c8",x"49",x"6b",x"7b"),
   130 => (x"71",x"b1",x"72",x"32"),
   131 => (x"26",x"4b",x"26",x"48"),
   132 => (x"5b",x"5e",x"0e",x"4f"),
   133 => (x"71",x"0e",x"5d",x"5c"),
   134 => (x"4c",x"d4",x"ff",x"4d"),
   135 => (x"ff",x"c3",x"48",x"75"),
   136 => (x"c2",x"7c",x"70",x"98"),
   137 => (x"05",x"bf",x"f4",x"e9"),
   138 => (x"66",x"d0",x"87",x"c8"),
   139 => (x"d4",x"30",x"c9",x"48"),
   140 => (x"66",x"d0",x"58",x"a6"),
   141 => (x"71",x"29",x"d8",x"49"),
   142 => (x"98",x"ff",x"c3",x"48"),
   143 => (x"66",x"d0",x"7c",x"70"),
   144 => (x"71",x"29",x"d0",x"49"),
   145 => (x"98",x"ff",x"c3",x"48"),
   146 => (x"66",x"d0",x"7c",x"70"),
   147 => (x"71",x"29",x"c8",x"49"),
   148 => (x"98",x"ff",x"c3",x"48"),
   149 => (x"66",x"d0",x"7c",x"70"),
   150 => (x"98",x"ff",x"c3",x"48"),
   151 => (x"49",x"75",x"7c",x"70"),
   152 => (x"48",x"71",x"29",x"d0"),
   153 => (x"70",x"98",x"ff",x"c3"),
   154 => (x"c9",x"4b",x"6c",x"7c"),
   155 => (x"c3",x"4a",x"ff",x"f0"),
   156 => (x"cf",x"05",x"ab",x"ff"),
   157 => (x"7c",x"71",x"49",x"87"),
   158 => (x"8a",x"c1",x"4b",x"6c"),
   159 => (x"71",x"87",x"c5",x"02"),
   160 => (x"87",x"f2",x"02",x"ab"),
   161 => (x"4d",x"26",x"48",x"73"),
   162 => (x"4b",x"26",x"4c",x"26"),
   163 => (x"c0",x"1e",x"4f",x"26"),
   164 => (x"48",x"d4",x"ff",x"49"),
   165 => (x"c1",x"78",x"ff",x"c3"),
   166 => (x"b7",x"c8",x"c3",x"81"),
   167 => (x"87",x"f1",x"04",x"a9"),
   168 => (x"5e",x"0e",x"4f",x"26"),
   169 => (x"0e",x"5d",x"5c",x"5b"),
   170 => (x"c1",x"f0",x"ff",x"c0"),
   171 => (x"c0",x"c1",x"4d",x"f7"),
   172 => (x"c0",x"c0",x"c0",x"c0"),
   173 => (x"87",x"d6",x"ff",x"4b"),
   174 => (x"4c",x"df",x"f8",x"c4"),
   175 => (x"49",x"75",x"1e",x"c0"),
   176 => (x"c4",x"87",x"ce",x"fd"),
   177 => (x"05",x"a8",x"c1",x"86"),
   178 => (x"ff",x"87",x"e5",x"c0"),
   179 => (x"ff",x"c3",x"48",x"d4"),
   180 => (x"c0",x"1e",x"73",x"78"),
   181 => (x"e9",x"c1",x"f0",x"e1"),
   182 => (x"87",x"f5",x"fc",x"49"),
   183 => (x"98",x"70",x"86",x"c4"),
   184 => (x"ff",x"87",x"ca",x"05"),
   185 => (x"ff",x"c3",x"48",x"d4"),
   186 => (x"cb",x"48",x"c1",x"78"),
   187 => (x"87",x"de",x"fe",x"87"),
   188 => (x"ff",x"05",x"8c",x"c1"),
   189 => (x"48",x"c0",x"87",x"c6"),
   190 => (x"4c",x"26",x"4d",x"26"),
   191 => (x"4f",x"26",x"4b",x"26"),
   192 => (x"5c",x"5b",x"5e",x"0e"),
   193 => (x"f0",x"ff",x"c0",x"0e"),
   194 => (x"ff",x"4c",x"c1",x"c1"),
   195 => (x"ff",x"c3",x"48",x"d4"),
   196 => (x"49",x"c4",x"cd",x"78"),
   197 => (x"d3",x"87",x"d0",x"f6"),
   198 => (x"74",x"1e",x"c0",x"4b"),
   199 => (x"87",x"f1",x"fb",x"49"),
   200 => (x"98",x"70",x"86",x"c4"),
   201 => (x"ff",x"87",x"ca",x"05"),
   202 => (x"ff",x"c3",x"48",x"d4"),
   203 => (x"cb",x"48",x"c1",x"78"),
   204 => (x"87",x"da",x"fd",x"87"),
   205 => (x"ff",x"05",x"8b",x"c1"),
   206 => (x"48",x"c0",x"87",x"df"),
   207 => (x"4b",x"26",x"4c",x"26"),
   208 => (x"00",x"00",x"4f",x"26"),
   209 => (x"00",x"44",x"4d",x"43"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"ff",x"c3",x"0e",x"5d"),
   212 => (x"4b",x"d4",x"ff",x"4d"),
   213 => (x"c6",x"87",x"f7",x"fc"),
   214 => (x"e1",x"c0",x"1e",x"ea"),
   215 => (x"49",x"c8",x"c1",x"f0"),
   216 => (x"c4",x"87",x"ee",x"fa"),
   217 => (x"02",x"a8",x"c1",x"86"),
   218 => (x"d3",x"fe",x"87",x"c8"),
   219 => (x"c1",x"48",x"c0",x"87"),
   220 => (x"f0",x"f9",x"87",x"e8"),
   221 => (x"cf",x"49",x"70",x"87"),
   222 => (x"c6",x"99",x"ff",x"ff"),
   223 => (x"c8",x"02",x"a9",x"ea"),
   224 => (x"87",x"fc",x"fd",x"87"),
   225 => (x"d1",x"c1",x"48",x"c0"),
   226 => (x"c0",x"7b",x"75",x"87"),
   227 => (x"d1",x"fc",x"4c",x"f1"),
   228 => (x"02",x"98",x"70",x"87"),
   229 => (x"c0",x"87",x"ec",x"c0"),
   230 => (x"f0",x"ff",x"c0",x"1e"),
   231 => (x"f9",x"49",x"fa",x"c1"),
   232 => (x"86",x"c4",x"87",x"ef"),
   233 => (x"da",x"05",x"98",x"70"),
   234 => (x"6b",x"7b",x"75",x"87"),
   235 => (x"75",x"7b",x"75",x"49"),
   236 => (x"75",x"7b",x"75",x"7b"),
   237 => (x"99",x"c0",x"c1",x"7b"),
   238 => (x"c1",x"87",x"c4",x"02"),
   239 => (x"c0",x"87",x"db",x"48"),
   240 => (x"c2",x"87",x"d7",x"48"),
   241 => (x"87",x"ca",x"05",x"ac"),
   242 => (x"f3",x"49",x"e4",x"cf"),
   243 => (x"48",x"c0",x"87",x"d9"),
   244 => (x"8c",x"c1",x"87",x"c8"),
   245 => (x"87",x"f6",x"fe",x"05"),
   246 => (x"4d",x"26",x"48",x"c0"),
   247 => (x"4b",x"26",x"4c",x"26"),
   248 => (x"00",x"00",x"4f",x"26"),
   249 => (x"43",x"48",x"44",x"53"),
   250 => (x"69",x"61",x"66",x"20"),
   251 => (x"00",x"0a",x"21",x"6c"),
   252 => (x"5c",x"5b",x"5e",x"0e"),
   253 => (x"d0",x"ff",x"0e",x"5d"),
   254 => (x"d0",x"e5",x"c0",x"4d"),
   255 => (x"c2",x"4c",x"c0",x"c1"),
   256 => (x"c1",x"48",x"f4",x"e9"),
   257 => (x"49",x"fc",x"d1",x"78"),
   258 => (x"c7",x"87",x"dc",x"f2"),
   259 => (x"f9",x"7d",x"c2",x"4b"),
   260 => (x"7d",x"c3",x"87",x"fc"),
   261 => (x"49",x"74",x"1e",x"c0"),
   262 => (x"c4",x"87",x"f6",x"f7"),
   263 => (x"05",x"a8",x"c1",x"86"),
   264 => (x"c2",x"4b",x"87",x"c1"),
   265 => (x"87",x"cb",x"05",x"ab"),
   266 => (x"f1",x"49",x"f4",x"d1"),
   267 => (x"48",x"c0",x"87",x"f9"),
   268 => (x"c1",x"87",x"f6",x"c0"),
   269 => (x"d4",x"ff",x"05",x"8b"),
   270 => (x"87",x"cc",x"fc",x"87"),
   271 => (x"58",x"f8",x"e9",x"c2"),
   272 => (x"cd",x"05",x"98",x"70"),
   273 => (x"c0",x"1e",x"c1",x"87"),
   274 => (x"d0",x"c1",x"f0",x"ff"),
   275 => (x"87",x"c1",x"f7",x"49"),
   276 => (x"d4",x"ff",x"86",x"c4"),
   277 => (x"78",x"ff",x"c3",x"48"),
   278 => (x"c2",x"87",x"cc",x"c5"),
   279 => (x"c2",x"58",x"fc",x"e9"),
   280 => (x"48",x"d4",x"ff",x"7d"),
   281 => (x"c1",x"78",x"ff",x"c3"),
   282 => (x"26",x"4d",x"26",x"48"),
   283 => (x"26",x"4b",x"26",x"4c"),
   284 => (x"00",x"00",x"00",x"4f"),
   285 => (x"52",x"52",x"45",x"49"),
   286 => (x"00",x"00",x"00",x"00"),
   287 => (x"00",x"49",x"50",x"53"),
   288 => (x"5c",x"5b",x"5e",x"0e"),
   289 => (x"4d",x"71",x"0e",x"5d"),
   290 => (x"ff",x"4c",x"ff",x"c3"),
   291 => (x"7b",x"74",x"4b",x"d4"),
   292 => (x"c4",x"48",x"d0",x"ff"),
   293 => (x"7b",x"74",x"78",x"c3"),
   294 => (x"ff",x"c0",x"1e",x"75"),
   295 => (x"49",x"d8",x"c1",x"f0"),
   296 => (x"c4",x"87",x"ee",x"f5"),
   297 => (x"02",x"98",x"70",x"86"),
   298 => (x"ec",x"d3",x"87",x"cb"),
   299 => (x"87",x"f7",x"ef",x"49"),
   300 => (x"ee",x"c0",x"48",x"c1"),
   301 => (x"c3",x"7b",x"74",x"87"),
   302 => (x"c0",x"c8",x"7b",x"fe"),
   303 => (x"49",x"66",x"d4",x"1e"),
   304 => (x"c4",x"87",x"d6",x"f3"),
   305 => (x"74",x"7b",x"74",x"86"),
   306 => (x"d8",x"7b",x"74",x"7b"),
   307 => (x"74",x"4a",x"e0",x"da"),
   308 => (x"c5",x"05",x"6b",x"7b"),
   309 => (x"05",x"8a",x"c1",x"87"),
   310 => (x"7b",x"74",x"87",x"f5"),
   311 => (x"c2",x"48",x"d0",x"ff"),
   312 => (x"26",x"48",x"c0",x"78"),
   313 => (x"26",x"4c",x"26",x"4d"),
   314 => (x"00",x"4f",x"26",x"4b"),
   315 => (x"74",x"69",x"72",x"57"),
   316 => (x"61",x"66",x"20",x"65"),
   317 => (x"64",x"65",x"6c",x"69"),
   318 => (x"5e",x"0e",x"00",x"0a"),
   319 => (x"0e",x"5d",x"5c",x"5b"),
   320 => (x"4b",x"71",x"86",x"fc"),
   321 => (x"c0",x"4c",x"d4",x"ff"),
   322 => (x"cd",x"ee",x"c5",x"7e"),
   323 => (x"ff",x"c3",x"4a",x"df"),
   324 => (x"c3",x"48",x"6c",x"7c"),
   325 => (x"c0",x"05",x"a8",x"fe"),
   326 => (x"4d",x"74",x"87",x"f8"),
   327 => (x"cc",x"02",x"9b",x"73"),
   328 => (x"1e",x"66",x"d4",x"87"),
   329 => (x"d3",x"f2",x"49",x"73"),
   330 => (x"d4",x"86",x"c4",x"87"),
   331 => (x"48",x"d0",x"ff",x"87"),
   332 => (x"d4",x"78",x"d1",x"c4"),
   333 => (x"ff",x"c3",x"4a",x"66"),
   334 => (x"05",x"8a",x"c1",x"7d"),
   335 => (x"a6",x"d8",x"87",x"f8"),
   336 => (x"7c",x"ff",x"c3",x"5a"),
   337 => (x"05",x"9b",x"73",x"7c"),
   338 => (x"d0",x"ff",x"87",x"c5"),
   339 => (x"c1",x"78",x"d0",x"48"),
   340 => (x"8a",x"c1",x"7e",x"4a"),
   341 => (x"87",x"f6",x"fe",x"05"),
   342 => (x"8e",x"fc",x"48",x"6e"),
   343 => (x"4c",x"26",x"4d",x"26"),
   344 => (x"4f",x"26",x"4b",x"26"),
   345 => (x"71",x"1e",x"73",x"1e"),
   346 => (x"ff",x"4b",x"c0",x"4a"),
   347 => (x"ff",x"c3",x"48",x"d4"),
   348 => (x"48",x"d0",x"ff",x"78"),
   349 => (x"ff",x"78",x"c3",x"c4"),
   350 => (x"ff",x"c3",x"48",x"d4"),
   351 => (x"c0",x"1e",x"72",x"78"),
   352 => (x"d1",x"c1",x"f0",x"ff"),
   353 => (x"87",x"c9",x"f2",x"49"),
   354 => (x"98",x"70",x"86",x"c4"),
   355 => (x"c8",x"87",x"d2",x"05"),
   356 => (x"66",x"cc",x"1e",x"c0"),
   357 => (x"87",x"e2",x"fd",x"49"),
   358 => (x"4b",x"70",x"86",x"c4"),
   359 => (x"c2",x"48",x"d0",x"ff"),
   360 => (x"26",x"48",x"73",x"78"),
   361 => (x"0e",x"4f",x"26",x"4b"),
   362 => (x"5d",x"5c",x"5b",x"5e"),
   363 => (x"c0",x"1e",x"c0",x"0e"),
   364 => (x"c9",x"c1",x"f0",x"ff"),
   365 => (x"87",x"d9",x"f1",x"49"),
   366 => (x"e9",x"c2",x"1e",x"d2"),
   367 => (x"f9",x"fc",x"49",x"fc"),
   368 => (x"c0",x"86",x"c8",x"87"),
   369 => (x"d2",x"84",x"c1",x"4c"),
   370 => (x"f8",x"04",x"ac",x"b7"),
   371 => (x"fc",x"e9",x"c2",x"87"),
   372 => (x"c3",x"49",x"bf",x"97"),
   373 => (x"c0",x"c1",x"99",x"c0"),
   374 => (x"e7",x"c0",x"05",x"a9"),
   375 => (x"c3",x"ea",x"c2",x"87"),
   376 => (x"d0",x"49",x"bf",x"97"),
   377 => (x"c4",x"ea",x"c2",x"31"),
   378 => (x"c8",x"4a",x"bf",x"97"),
   379 => (x"c2",x"b1",x"72",x"32"),
   380 => (x"bf",x"97",x"c5",x"ea"),
   381 => (x"4c",x"71",x"b1",x"4a"),
   382 => (x"ff",x"ff",x"ff",x"cf"),
   383 => (x"ca",x"84",x"c1",x"9c"),
   384 => (x"87",x"e7",x"c1",x"34"),
   385 => (x"97",x"c5",x"ea",x"c2"),
   386 => (x"31",x"c1",x"49",x"bf"),
   387 => (x"ea",x"c2",x"99",x"c6"),
   388 => (x"4a",x"bf",x"97",x"c6"),
   389 => (x"72",x"2a",x"b7",x"c7"),
   390 => (x"c1",x"ea",x"c2",x"b1"),
   391 => (x"4d",x"4a",x"bf",x"97"),
   392 => (x"ea",x"c2",x"9d",x"cf"),
   393 => (x"4a",x"bf",x"97",x"c2"),
   394 => (x"32",x"ca",x"9a",x"c3"),
   395 => (x"97",x"c3",x"ea",x"c2"),
   396 => (x"33",x"c2",x"4b",x"bf"),
   397 => (x"ea",x"c2",x"b2",x"73"),
   398 => (x"4b",x"bf",x"97",x"c4"),
   399 => (x"c6",x"9b",x"c0",x"c3"),
   400 => (x"b2",x"73",x"2b",x"b7"),
   401 => (x"48",x"c1",x"81",x"c2"),
   402 => (x"49",x"70",x"30",x"71"),
   403 => (x"30",x"75",x"48",x"c1"),
   404 => (x"4c",x"72",x"4d",x"70"),
   405 => (x"94",x"71",x"84",x"c1"),
   406 => (x"ad",x"b7",x"c0",x"c8"),
   407 => (x"c1",x"87",x"cc",x"06"),
   408 => (x"c8",x"2d",x"b7",x"34"),
   409 => (x"01",x"ad",x"b7",x"c0"),
   410 => (x"74",x"87",x"f4",x"ff"),
   411 => (x"26",x"4d",x"26",x"48"),
   412 => (x"26",x"4b",x"26",x"4c"),
   413 => (x"5b",x"5e",x"0e",x"4f"),
   414 => (x"f8",x"0e",x"5d",x"5c"),
   415 => (x"e4",x"f2",x"c2",x"86"),
   416 => (x"c2",x"78",x"c0",x"48"),
   417 => (x"c0",x"1e",x"dc",x"ea"),
   418 => (x"87",x"d8",x"fb",x"49"),
   419 => (x"98",x"70",x"86",x"c4"),
   420 => (x"c0",x"87",x"c5",x"05"),
   421 => (x"87",x"c0",x"c9",x"48"),
   422 => (x"7e",x"c1",x"4d",x"c0"),
   423 => (x"bf",x"c0",x"ff",x"c0"),
   424 => (x"d2",x"eb",x"c2",x"49"),
   425 => (x"4b",x"c8",x"71",x"4a"),
   426 => (x"70",x"87",x"fb",x"e8"),
   427 => (x"87",x"c2",x"05",x"98"),
   428 => (x"fe",x"c0",x"7e",x"c0"),
   429 => (x"c2",x"49",x"bf",x"fc"),
   430 => (x"71",x"4a",x"ee",x"eb"),
   431 => (x"e5",x"e8",x"4b",x"c8"),
   432 => (x"05",x"98",x"70",x"87"),
   433 => (x"7e",x"c0",x"87",x"c2"),
   434 => (x"fd",x"c0",x"02",x"6e"),
   435 => (x"e2",x"f1",x"c2",x"87"),
   436 => (x"f2",x"c2",x"4d",x"bf"),
   437 => (x"7e",x"bf",x"9f",x"da"),
   438 => (x"ea",x"d6",x"c5",x"48"),
   439 => (x"87",x"c7",x"05",x"a8"),
   440 => (x"bf",x"e2",x"f1",x"c2"),
   441 => (x"6e",x"87",x"ce",x"4d"),
   442 => (x"d5",x"e9",x"ca",x"48"),
   443 => (x"87",x"c5",x"02",x"a8"),
   444 => (x"e3",x"c7",x"48",x"c0"),
   445 => (x"dc",x"ea",x"c2",x"87"),
   446 => (x"f9",x"49",x"75",x"1e"),
   447 => (x"86",x"c4",x"87",x"e6"),
   448 => (x"c5",x"05",x"98",x"70"),
   449 => (x"c7",x"48",x"c0",x"87"),
   450 => (x"fe",x"c0",x"87",x"ce"),
   451 => (x"c2",x"49",x"bf",x"fc"),
   452 => (x"71",x"4a",x"ee",x"eb"),
   453 => (x"cd",x"e7",x"4b",x"c8"),
   454 => (x"05",x"98",x"70",x"87"),
   455 => (x"f2",x"c2",x"87",x"c8"),
   456 => (x"78",x"c1",x"48",x"e4"),
   457 => (x"ff",x"c0",x"87",x"da"),
   458 => (x"c2",x"49",x"bf",x"c0"),
   459 => (x"71",x"4a",x"d2",x"eb"),
   460 => (x"f1",x"e6",x"4b",x"c8"),
   461 => (x"02",x"98",x"70",x"87"),
   462 => (x"c0",x"87",x"c5",x"c0"),
   463 => (x"87",x"d8",x"c6",x"48"),
   464 => (x"97",x"da",x"f2",x"c2"),
   465 => (x"d5",x"c1",x"49",x"bf"),
   466 => (x"cd",x"c0",x"05",x"a9"),
   467 => (x"db",x"f2",x"c2",x"87"),
   468 => (x"c2",x"49",x"bf",x"97"),
   469 => (x"c0",x"02",x"a9",x"ea"),
   470 => (x"48",x"c0",x"87",x"c5"),
   471 => (x"c2",x"87",x"f9",x"c5"),
   472 => (x"bf",x"97",x"dc",x"ea"),
   473 => (x"e9",x"c3",x"48",x"7e"),
   474 => (x"ce",x"c0",x"02",x"a8"),
   475 => (x"c3",x"48",x"6e",x"87"),
   476 => (x"c0",x"02",x"a8",x"eb"),
   477 => (x"48",x"c0",x"87",x"c5"),
   478 => (x"c2",x"87",x"dd",x"c5"),
   479 => (x"bf",x"97",x"e7",x"ea"),
   480 => (x"c0",x"05",x"99",x"49"),
   481 => (x"ea",x"c2",x"87",x"cc"),
   482 => (x"49",x"bf",x"97",x"e8"),
   483 => (x"c0",x"02",x"a9",x"c2"),
   484 => (x"48",x"c0",x"87",x"c5"),
   485 => (x"c2",x"87",x"c1",x"c5"),
   486 => (x"bf",x"97",x"e9",x"ea"),
   487 => (x"e0",x"f2",x"c2",x"48"),
   488 => (x"48",x"4c",x"70",x"58"),
   489 => (x"f2",x"c2",x"88",x"c1"),
   490 => (x"ea",x"c2",x"58",x"e4"),
   491 => (x"49",x"bf",x"97",x"ea"),
   492 => (x"ea",x"c2",x"81",x"75"),
   493 => (x"4a",x"bf",x"97",x"eb"),
   494 => (x"a1",x"72",x"32",x"c8"),
   495 => (x"f4",x"f6",x"c2",x"7e"),
   496 => (x"c2",x"78",x"6e",x"48"),
   497 => (x"bf",x"97",x"ec",x"ea"),
   498 => (x"58",x"a6",x"c8",x"48"),
   499 => (x"bf",x"e4",x"f2",x"c2"),
   500 => (x"87",x"cf",x"c2",x"02"),
   501 => (x"bf",x"fc",x"fe",x"c0"),
   502 => (x"ee",x"eb",x"c2",x"49"),
   503 => (x"4b",x"c8",x"71",x"4a"),
   504 => (x"70",x"87",x"c3",x"e4"),
   505 => (x"c5",x"c0",x"02",x"98"),
   506 => (x"c3",x"48",x"c0",x"87"),
   507 => (x"f2",x"c2",x"87",x"ea"),
   508 => (x"c2",x"4c",x"bf",x"dc"),
   509 => (x"c2",x"5c",x"c8",x"f7"),
   510 => (x"bf",x"97",x"c1",x"eb"),
   511 => (x"c2",x"31",x"c8",x"49"),
   512 => (x"bf",x"97",x"c0",x"eb"),
   513 => (x"c2",x"49",x"a1",x"4a"),
   514 => (x"bf",x"97",x"c2",x"eb"),
   515 => (x"72",x"32",x"d0",x"4a"),
   516 => (x"eb",x"c2",x"49",x"a1"),
   517 => (x"4a",x"bf",x"97",x"c3"),
   518 => (x"a1",x"72",x"32",x"d8"),
   519 => (x"91",x"66",x"c4",x"49"),
   520 => (x"bf",x"f4",x"f6",x"c2"),
   521 => (x"fc",x"f6",x"c2",x"81"),
   522 => (x"c9",x"eb",x"c2",x"59"),
   523 => (x"c8",x"4a",x"bf",x"97"),
   524 => (x"c8",x"eb",x"c2",x"32"),
   525 => (x"a2",x"4b",x"bf",x"97"),
   526 => (x"ca",x"eb",x"c2",x"4a"),
   527 => (x"d0",x"4b",x"bf",x"97"),
   528 => (x"4a",x"a2",x"73",x"33"),
   529 => (x"97",x"cb",x"eb",x"c2"),
   530 => (x"9b",x"cf",x"4b",x"bf"),
   531 => (x"a2",x"73",x"33",x"d8"),
   532 => (x"c0",x"f7",x"c2",x"4a"),
   533 => (x"74",x"8a",x"c2",x"5a"),
   534 => (x"c0",x"f7",x"c2",x"92"),
   535 => (x"78",x"a1",x"72",x"48"),
   536 => (x"c2",x"87",x"c1",x"c1"),
   537 => (x"bf",x"97",x"ee",x"ea"),
   538 => (x"c2",x"31",x"c8",x"49"),
   539 => (x"bf",x"97",x"ed",x"ea"),
   540 => (x"c5",x"49",x"a1",x"4a"),
   541 => (x"81",x"ff",x"c7",x"31"),
   542 => (x"f7",x"c2",x"29",x"c9"),
   543 => (x"ea",x"c2",x"59",x"c8"),
   544 => (x"4a",x"bf",x"97",x"f3"),
   545 => (x"ea",x"c2",x"32",x"c8"),
   546 => (x"4b",x"bf",x"97",x"f2"),
   547 => (x"66",x"c4",x"4a",x"a2"),
   548 => (x"c2",x"82",x"6e",x"92"),
   549 => (x"c2",x"5a",x"c4",x"f7"),
   550 => (x"c0",x"48",x"fc",x"f6"),
   551 => (x"f8",x"f6",x"c2",x"78"),
   552 => (x"78",x"a1",x"72",x"48"),
   553 => (x"48",x"c8",x"f7",x"c2"),
   554 => (x"bf",x"fc",x"f6",x"c2"),
   555 => (x"cc",x"f7",x"c2",x"78"),
   556 => (x"c0",x"f7",x"c2",x"48"),
   557 => (x"f2",x"c2",x"78",x"bf"),
   558 => (x"c0",x"02",x"bf",x"e4"),
   559 => (x"48",x"74",x"87",x"c9"),
   560 => (x"7e",x"70",x"30",x"c4"),
   561 => (x"c2",x"87",x"c9",x"c0"),
   562 => (x"48",x"bf",x"c4",x"f7"),
   563 => (x"7e",x"70",x"30",x"c4"),
   564 => (x"48",x"e8",x"f2",x"c2"),
   565 => (x"48",x"c1",x"78",x"6e"),
   566 => (x"4d",x"26",x"8e",x"f8"),
   567 => (x"4b",x"26",x"4c",x"26"),
   568 => (x"5e",x"0e",x"4f",x"26"),
   569 => (x"0e",x"5d",x"5c",x"5b"),
   570 => (x"f2",x"c2",x"4a",x"71"),
   571 => (x"cb",x"02",x"bf",x"e4"),
   572 => (x"c7",x"4b",x"72",x"87"),
   573 => (x"c1",x"4d",x"72",x"2b"),
   574 => (x"87",x"c9",x"9d",x"ff"),
   575 => (x"2b",x"c8",x"4b",x"72"),
   576 => (x"ff",x"c3",x"4d",x"72"),
   577 => (x"f4",x"f6",x"c2",x"9d"),
   578 => (x"fe",x"c0",x"83",x"bf"),
   579 => (x"02",x"ab",x"bf",x"f8"),
   580 => (x"fe",x"c0",x"87",x"d9"),
   581 => (x"ea",x"c2",x"5b",x"fc"),
   582 => (x"49",x"73",x"1e",x"dc"),
   583 => (x"c4",x"87",x"c5",x"f1"),
   584 => (x"05",x"98",x"70",x"86"),
   585 => (x"48",x"c0",x"87",x"c5"),
   586 => (x"c2",x"87",x"e6",x"c0"),
   587 => (x"02",x"bf",x"e4",x"f2"),
   588 => (x"49",x"75",x"87",x"d2"),
   589 => (x"ea",x"c2",x"91",x"c4"),
   590 => (x"4c",x"69",x"81",x"dc"),
   591 => (x"ff",x"ff",x"ff",x"cf"),
   592 => (x"87",x"cb",x"9c",x"ff"),
   593 => (x"91",x"c2",x"49",x"75"),
   594 => (x"81",x"dc",x"ea",x"c2"),
   595 => (x"74",x"4c",x"69",x"9f"),
   596 => (x"26",x"4d",x"26",x"48"),
   597 => (x"26",x"4b",x"26",x"4c"),
   598 => (x"5b",x"5e",x"0e",x"4f"),
   599 => (x"f0",x"0e",x"5d",x"5c"),
   600 => (x"59",x"a6",x"cc",x"86"),
   601 => (x"c5",x"05",x"66",x"c8"),
   602 => (x"c4",x"48",x"c0",x"87"),
   603 => (x"66",x"c8",x"87",x"c4"),
   604 => (x"70",x"80",x"c8",x"48"),
   605 => (x"78",x"c0",x"48",x"7e"),
   606 => (x"02",x"66",x"e0",x"c0"),
   607 => (x"e0",x"c0",x"87",x"c8"),
   608 => (x"05",x"bf",x"97",x"66"),
   609 => (x"48",x"c0",x"87",x"c5"),
   610 => (x"c0",x"87",x"e7",x"c3"),
   611 => (x"49",x"49",x"c1",x"1e"),
   612 => (x"c4",x"87",x"ea",x"d0"),
   613 => (x"9c",x"4c",x"70",x"86"),
   614 => (x"87",x"fe",x"c0",x"02"),
   615 => (x"4a",x"ec",x"f2",x"c2"),
   616 => (x"49",x"66",x"e0",x"c0"),
   617 => (x"87",x"e3",x"dc",x"ff"),
   618 => (x"c0",x"02",x"98",x"70"),
   619 => (x"4a",x"74",x"87",x"ec"),
   620 => (x"49",x"66",x"e0",x"c0"),
   621 => (x"dd",x"ff",x"4b",x"cb"),
   622 => (x"98",x"70",x"87",x"c6"),
   623 => (x"c0",x"87",x"db",x"02"),
   624 => (x"02",x"9c",x"74",x"1e"),
   625 => (x"4d",x"c0",x"87",x"c4"),
   626 => (x"4d",x"c1",x"87",x"c2"),
   627 => (x"ec",x"cf",x"49",x"75"),
   628 => (x"70",x"86",x"c4",x"87"),
   629 => (x"ff",x"05",x"9c",x"4c"),
   630 => (x"9c",x"74",x"87",x"c2"),
   631 => (x"87",x"d0",x"c2",x"02"),
   632 => (x"6e",x"49",x"a4",x"dc"),
   633 => (x"da",x"78",x"69",x"48"),
   634 => (x"66",x"c8",x"49",x"a4"),
   635 => (x"c8",x"80",x"c4",x"48"),
   636 => (x"69",x"9f",x"58",x"a6"),
   637 => (x"08",x"66",x"c4",x"48"),
   638 => (x"e4",x"f2",x"c2",x"78"),
   639 => (x"87",x"d2",x"02",x"bf"),
   640 => (x"9f",x"49",x"a4",x"d4"),
   641 => (x"ff",x"c0",x"49",x"69"),
   642 => (x"48",x"71",x"99",x"ff"),
   643 => (x"58",x"a6",x"30",x"d0"),
   644 => (x"a6",x"cc",x"87",x"c5"),
   645 => (x"cc",x"78",x"c0",x"48"),
   646 => (x"66",x"c4",x"48",x"66"),
   647 => (x"66",x"c4",x"80",x"bf"),
   648 => (x"66",x"c8",x"78",x"08"),
   649 => (x"c8",x"78",x"c0",x"48"),
   650 => (x"81",x"cc",x"49",x"66"),
   651 => (x"79",x"bf",x"66",x"c4"),
   652 => (x"d0",x"49",x"66",x"c8"),
   653 => (x"4d",x"79",x"c0",x"81"),
   654 => (x"c8",x"4c",x"66",x"c4"),
   655 => (x"82",x"d4",x"4a",x"66"),
   656 => (x"91",x"c8",x"49",x"75"),
   657 => (x"c0",x"49",x"a1",x"72"),
   658 => (x"c1",x"79",x"6c",x"41"),
   659 => (x"ad",x"b7",x"c6",x"85"),
   660 => (x"87",x"e7",x"ff",x"04"),
   661 => (x"c9",x"4a",x"bf",x"6e"),
   662 => (x"c0",x"49",x"72",x"2a"),
   663 => (x"db",x"ff",x"4a",x"f0"),
   664 => (x"4a",x"70",x"87",x"d2"),
   665 => (x"c1",x"49",x"66",x"c8"),
   666 => (x"79",x"72",x"81",x"c4"),
   667 => (x"87",x"c2",x"48",x"c1"),
   668 => (x"8e",x"f0",x"48",x"c0"),
   669 => (x"4c",x"26",x"4d",x"26"),
   670 => (x"4f",x"26",x"4b",x"26"),
   671 => (x"5c",x"5b",x"5e",x"0e"),
   672 => (x"4c",x"71",x"0e",x"5d"),
   673 => (x"74",x"4d",x"66",x"d0"),
   674 => (x"c2",x"c1",x"02",x"9c"),
   675 => (x"49",x"a4",x"c8",x"87"),
   676 => (x"fa",x"c0",x"02",x"69"),
   677 => (x"85",x"49",x"6c",x"87"),
   678 => (x"f2",x"c2",x"b9",x"75"),
   679 => (x"ff",x"4a",x"bf",x"e0"),
   680 => (x"71",x"99",x"72",x"ba"),
   681 => (x"e4",x"c0",x"02",x"99"),
   682 => (x"4b",x"a4",x"c4",x"87"),
   683 => (x"f1",x"f8",x"49",x"6b"),
   684 => (x"c2",x"7b",x"70",x"87"),
   685 => (x"49",x"bf",x"dc",x"f2"),
   686 => (x"7c",x"71",x"81",x"6c"),
   687 => (x"f2",x"c2",x"b9",x"75"),
   688 => (x"ff",x"4a",x"bf",x"e0"),
   689 => (x"71",x"99",x"72",x"ba"),
   690 => (x"dc",x"ff",x"05",x"99"),
   691 => (x"26",x"7c",x"75",x"87"),
   692 => (x"26",x"4c",x"26",x"4d"),
   693 => (x"1e",x"4f",x"26",x"4b"),
   694 => (x"4b",x"71",x"1e",x"73"),
   695 => (x"87",x"c7",x"02",x"9b"),
   696 => (x"69",x"49",x"a3",x"c8"),
   697 => (x"c0",x"87",x"c5",x"05"),
   698 => (x"87",x"f6",x"c0",x"48"),
   699 => (x"bf",x"f8",x"f6",x"c2"),
   700 => (x"4a",x"a3",x"c4",x"49"),
   701 => (x"8a",x"c2",x"4a",x"6a"),
   702 => (x"bf",x"dc",x"f2",x"c2"),
   703 => (x"49",x"a1",x"72",x"92"),
   704 => (x"bf",x"e0",x"f2",x"c2"),
   705 => (x"72",x"9a",x"6b",x"4a"),
   706 => (x"fe",x"c0",x"49",x"a1"),
   707 => (x"66",x"c8",x"59",x"fc"),
   708 => (x"cf",x"e9",x"71",x"1e"),
   709 => (x"70",x"86",x"c4",x"87"),
   710 => (x"87",x"c4",x"05",x"98"),
   711 => (x"87",x"c2",x"48",x"c0"),
   712 => (x"4b",x"26",x"48",x"c1"),
   713 => (x"73",x"1e",x"4f",x"26"),
   714 => (x"9b",x"4b",x"71",x"1e"),
   715 => (x"c8",x"87",x"c7",x"02"),
   716 => (x"05",x"69",x"49",x"a3"),
   717 => (x"48",x"c0",x"87",x"c5"),
   718 => (x"c2",x"87",x"f6",x"c0"),
   719 => (x"49",x"bf",x"f8",x"f6"),
   720 => (x"6a",x"4a",x"a3",x"c4"),
   721 => (x"c2",x"8a",x"c2",x"4a"),
   722 => (x"92",x"bf",x"dc",x"f2"),
   723 => (x"c2",x"49",x"a1",x"72"),
   724 => (x"4a",x"bf",x"e0",x"f2"),
   725 => (x"a1",x"72",x"9a",x"6b"),
   726 => (x"fc",x"fe",x"c0",x"49"),
   727 => (x"1e",x"66",x"c8",x"59"),
   728 => (x"87",x"dc",x"e4",x"71"),
   729 => (x"98",x"70",x"86",x"c4"),
   730 => (x"c0",x"87",x"c4",x"05"),
   731 => (x"c1",x"87",x"c2",x"48"),
   732 => (x"26",x"4b",x"26",x"48"),
   733 => (x"5b",x"5e",x"0e",x"4f"),
   734 => (x"f8",x"0e",x"5d",x"5c"),
   735 => (x"c4",x"7e",x"71",x"86"),
   736 => (x"78",x"ff",x"48",x"a6"),
   737 => (x"ff",x"ff",x"ff",x"c1"),
   738 => (x"c0",x"4d",x"ff",x"ff"),
   739 => (x"d4",x"4a",x"6e",x"4b"),
   740 => (x"c8",x"49",x"73",x"82"),
   741 => (x"49",x"a1",x"72",x"91"),
   742 => (x"69",x"4c",x"66",x"d8"),
   743 => (x"ac",x"b7",x"c0",x"8c"),
   744 => (x"75",x"87",x"cb",x"04"),
   745 => (x"c5",x"03",x"ac",x"b7"),
   746 => (x"5b",x"a6",x"c8",x"87"),
   747 => (x"83",x"c1",x"4d",x"74"),
   748 => (x"04",x"ab",x"b7",x"c6"),
   749 => (x"c4",x"87",x"d6",x"ff"),
   750 => (x"8e",x"f8",x"48",x"66"),
   751 => (x"4c",x"26",x"4d",x"26"),
   752 => (x"4f",x"26",x"4b",x"26"),
   753 => (x"5c",x"5b",x"5e",x"0e"),
   754 => (x"86",x"f0",x"0e",x"5d"),
   755 => (x"a6",x"c4",x"7e",x"71"),
   756 => (x"ff",x"ff",x"c1",x"48"),
   757 => (x"78",x"ff",x"ff",x"ff"),
   758 => (x"78",x"ff",x"80",x"c4"),
   759 => (x"4c",x"c0",x"4d",x"c0"),
   760 => (x"83",x"d4",x"4b",x"6e"),
   761 => (x"92",x"c8",x"4a",x"74"),
   762 => (x"75",x"4a",x"a2",x"73"),
   763 => (x"73",x"91",x"c8",x"49"),
   764 => (x"48",x"6a",x"49",x"a1"),
   765 => (x"49",x"70",x"88",x"69"),
   766 => (x"74",x"59",x"a6",x"d0"),
   767 => (x"87",x"d2",x"02",x"ad"),
   768 => (x"c4",x"48",x"66",x"cc"),
   769 => (x"c9",x"03",x"a8",x"66"),
   770 => (x"5c",x"a6",x"cc",x"87"),
   771 => (x"cc",x"48",x"a6",x"c4"),
   772 => (x"84",x"c1",x"78",x"66"),
   773 => (x"04",x"ac",x"b7",x"c6"),
   774 => (x"c1",x"87",x"c5",x"ff"),
   775 => (x"ad",x"b7",x"c6",x"85"),
   776 => (x"87",x"fa",x"fe",x"04"),
   777 => (x"f0",x"48",x"66",x"c8"),
   778 => (x"26",x"4d",x"26",x"8e"),
   779 => (x"26",x"4b",x"26",x"4c"),
   780 => (x"5b",x"5e",x"0e",x"4f"),
   781 => (x"ec",x"0e",x"5d",x"5c"),
   782 => (x"c0",x"4b",x"71",x"86"),
   783 => (x"c9",x"48",x"66",x"e4"),
   784 => (x"58",x"a6",x"c8",x"28"),
   785 => (x"bf",x"e0",x"f2",x"c2"),
   786 => (x"72",x"ba",x"ff",x"4a"),
   787 => (x"98",x"66",x"c4",x"48"),
   788 => (x"73",x"58",x"a6",x"cc"),
   789 => (x"c1",x"c3",x"02",x"9b"),
   790 => (x"49",x"a3",x"c8",x"87"),
   791 => (x"f9",x"c2",x"02",x"69"),
   792 => (x"6b",x"48",x"72",x"87"),
   793 => (x"58",x"a6",x"d4",x"98"),
   794 => (x"6c",x"4c",x"a3",x"c4"),
   795 => (x"48",x"66",x"c8",x"7e"),
   796 => (x"05",x"a8",x"66",x"d0"),
   797 => (x"66",x"c4",x"87",x"c6"),
   798 => (x"87",x"cc",x"c2",x"7b"),
   799 => (x"73",x"1e",x"66",x"c8"),
   800 => (x"87",x"f1",x"fb",x"49"),
   801 => (x"4d",x"70",x"86",x"c4"),
   802 => (x"04",x"ad",x"b7",x"c0"),
   803 => (x"a3",x"d4",x"87",x"d0"),
   804 => (x"c8",x"49",x"75",x"4a"),
   805 => (x"49",x"a1",x"72",x"91"),
   806 => (x"7c",x"69",x"7b",x"21"),
   807 => (x"7b",x"c0",x"87",x"c7"),
   808 => (x"69",x"49",x"a3",x"cc"),
   809 => (x"48",x"66",x"c4",x"7c"),
   810 => (x"a6",x"c8",x"88",x"6b"),
   811 => (x"1e",x"66",x"d0",x"58"),
   812 => (x"c0",x"fb",x"49",x"73"),
   813 => (x"70",x"86",x"c4",x"87"),
   814 => (x"a3",x"c4",x"c1",x"4d"),
   815 => (x"48",x"a6",x"c8",x"49"),
   816 => (x"66",x"d0",x"78",x"69"),
   817 => (x"a8",x"66",x"c8",x"48"),
   818 => (x"87",x"f2",x"c0",x"06"),
   819 => (x"04",x"ad",x"b7",x"c0"),
   820 => (x"cc",x"87",x"eb",x"c0"),
   821 => (x"a3",x"d4",x"48",x"a6"),
   822 => (x"c8",x"49",x"75",x"78"),
   823 => (x"81",x"66",x"cc",x"91"),
   824 => (x"69",x"48",x"66",x"d0"),
   825 => (x"c8",x"49",x"70",x"88"),
   826 => (x"d1",x"06",x"a9",x"66"),
   827 => (x"fb",x"49",x"73",x"87"),
   828 => (x"49",x"70",x"87",x"d2"),
   829 => (x"66",x"cc",x"91",x"c8"),
   830 => (x"41",x"66",x"d0",x"81"),
   831 => (x"66",x"c4",x"79",x"6e"),
   832 => (x"f5",x"49",x"73",x"1e"),
   833 => (x"86",x"c4",x"87",x"f6"),
   834 => (x"1e",x"dc",x"ea",x"c2"),
   835 => (x"c6",x"f7",x"49",x"73"),
   836 => (x"d0",x"86",x"c4",x"87"),
   837 => (x"e4",x"c0",x"49",x"a3"),
   838 => (x"8e",x"ec",x"79",x"66"),
   839 => (x"4c",x"26",x"4d",x"26"),
   840 => (x"4f",x"26",x"4b",x"26"),
   841 => (x"71",x"1e",x"73",x"1e"),
   842 => (x"c0",x"02",x"9b",x"4b"),
   843 => (x"f7",x"c2",x"87",x"e4"),
   844 => (x"4a",x"73",x"5b",x"cc"),
   845 => (x"f2",x"c2",x"8a",x"c2"),
   846 => (x"92",x"49",x"bf",x"dc"),
   847 => (x"bf",x"f8",x"f6",x"c2"),
   848 => (x"c2",x"80",x"72",x"48"),
   849 => (x"71",x"58",x"d0",x"f7"),
   850 => (x"c2",x"30",x"c4",x"48"),
   851 => (x"c0",x"58",x"ec",x"f2"),
   852 => (x"f7",x"c2",x"87",x"ed"),
   853 => (x"f6",x"c2",x"48",x"c8"),
   854 => (x"c2",x"78",x"bf",x"fc"),
   855 => (x"c2",x"48",x"cc",x"f7"),
   856 => (x"78",x"bf",x"c0",x"f7"),
   857 => (x"bf",x"e4",x"f2",x"c2"),
   858 => (x"c2",x"87",x"c9",x"02"),
   859 => (x"49",x"bf",x"dc",x"f2"),
   860 => (x"87",x"c7",x"31",x"c4"),
   861 => (x"bf",x"c4",x"f7",x"c2"),
   862 => (x"c2",x"31",x"c4",x"49"),
   863 => (x"26",x"59",x"ec",x"f2"),
   864 => (x"0e",x"4f",x"26",x"4b"),
   865 => (x"0e",x"5c",x"5b",x"5e"),
   866 => (x"4b",x"c0",x"4a",x"71"),
   867 => (x"c0",x"02",x"9a",x"72"),
   868 => (x"a2",x"da",x"87",x"e0"),
   869 => (x"4b",x"69",x"9f",x"49"),
   870 => (x"bf",x"e4",x"f2",x"c2"),
   871 => (x"d4",x"87",x"cf",x"02"),
   872 => (x"69",x"9f",x"49",x"a2"),
   873 => (x"ff",x"c0",x"4c",x"49"),
   874 => (x"34",x"d0",x"9c",x"ff"),
   875 => (x"4c",x"c0",x"87",x"c2"),
   876 => (x"49",x"73",x"b3",x"74"),
   877 => (x"26",x"87",x"ed",x"fd"),
   878 => (x"26",x"4b",x"26",x"4c"),
   879 => (x"5b",x"5e",x"0e",x"4f"),
   880 => (x"f0",x"0e",x"5d",x"5c"),
   881 => (x"59",x"a6",x"c8",x"86"),
   882 => (x"ff",x"ff",x"ff",x"cf"),
   883 => (x"7e",x"c0",x"4c",x"f8"),
   884 => (x"d8",x"02",x"66",x"c4"),
   885 => (x"d8",x"ea",x"c2",x"87"),
   886 => (x"c2",x"78",x"c0",x"48"),
   887 => (x"c2",x"48",x"d0",x"ea"),
   888 => (x"78",x"bf",x"cc",x"f7"),
   889 => (x"48",x"d4",x"ea",x"c2"),
   890 => (x"bf",x"c8",x"f7",x"c2"),
   891 => (x"f9",x"f2",x"c2",x"78"),
   892 => (x"c2",x"50",x"c0",x"48"),
   893 => (x"49",x"bf",x"e8",x"f2"),
   894 => (x"bf",x"d8",x"ea",x"c2"),
   895 => (x"03",x"aa",x"71",x"4a"),
   896 => (x"72",x"87",x"cc",x"c4"),
   897 => (x"05",x"99",x"cf",x"49"),
   898 => (x"c0",x"87",x"ea",x"c0"),
   899 => (x"c2",x"48",x"f8",x"fe"),
   900 => (x"78",x"bf",x"d0",x"ea"),
   901 => (x"1e",x"dc",x"ea",x"c2"),
   902 => (x"bf",x"d0",x"ea",x"c2"),
   903 => (x"d0",x"ea",x"c2",x"49"),
   904 => (x"78",x"a1",x"c1",x"48"),
   905 => (x"fb",x"dc",x"ff",x"71"),
   906 => (x"c0",x"86",x"c4",x"87"),
   907 => (x"c2",x"48",x"f4",x"fe"),
   908 => (x"cc",x"78",x"dc",x"ea"),
   909 => (x"f4",x"fe",x"c0",x"87"),
   910 => (x"e0",x"c0",x"48",x"bf"),
   911 => (x"f8",x"fe",x"c0",x"80"),
   912 => (x"d8",x"ea",x"c2",x"58"),
   913 => (x"80",x"c1",x"48",x"bf"),
   914 => (x"58",x"dc",x"ea",x"c2"),
   915 => (x"00",x"0f",x"b4",x"27"),
   916 => (x"bf",x"97",x"bf",x"00"),
   917 => (x"c2",x"02",x"9d",x"4d"),
   918 => (x"e5",x"c3",x"87",x"e5"),
   919 => (x"de",x"c2",x"02",x"ad"),
   920 => (x"f4",x"fe",x"c0",x"87"),
   921 => (x"a3",x"cb",x"4b",x"bf"),
   922 => (x"cf",x"4c",x"11",x"49"),
   923 => (x"d2",x"c1",x"05",x"ac"),
   924 => (x"df",x"49",x"75",x"87"),
   925 => (x"cd",x"89",x"c1",x"99"),
   926 => (x"ec",x"f2",x"c2",x"91"),
   927 => (x"4a",x"a3",x"c1",x"81"),
   928 => (x"a3",x"c3",x"51",x"12"),
   929 => (x"c5",x"51",x"12",x"4a"),
   930 => (x"51",x"12",x"4a",x"a3"),
   931 => (x"12",x"4a",x"a3",x"c7"),
   932 => (x"4a",x"a3",x"c9",x"51"),
   933 => (x"a3",x"ce",x"51",x"12"),
   934 => (x"d0",x"51",x"12",x"4a"),
   935 => (x"51",x"12",x"4a",x"a3"),
   936 => (x"12",x"4a",x"a3",x"d2"),
   937 => (x"4a",x"a3",x"d4",x"51"),
   938 => (x"a3",x"d6",x"51",x"12"),
   939 => (x"d8",x"51",x"12",x"4a"),
   940 => (x"51",x"12",x"4a",x"a3"),
   941 => (x"12",x"4a",x"a3",x"dc"),
   942 => (x"4a",x"a3",x"de",x"51"),
   943 => (x"7e",x"c1",x"51",x"12"),
   944 => (x"74",x"87",x"fc",x"c0"),
   945 => (x"05",x"99",x"c8",x"49"),
   946 => (x"74",x"87",x"ed",x"c0"),
   947 => (x"05",x"99",x"d0",x"49"),
   948 => (x"e0",x"c0",x"87",x"d3"),
   949 => (x"cc",x"c0",x"02",x"66"),
   950 => (x"c0",x"49",x"73",x"87"),
   951 => (x"70",x"0f",x"66",x"e0"),
   952 => (x"d3",x"c0",x"02",x"98"),
   953 => (x"c0",x"05",x"6e",x"87"),
   954 => (x"f2",x"c2",x"87",x"c6"),
   955 => (x"50",x"c0",x"48",x"ec"),
   956 => (x"bf",x"f4",x"fe",x"c0"),
   957 => (x"87",x"e9",x"c2",x"48"),
   958 => (x"48",x"f9",x"f2",x"c2"),
   959 => (x"c2",x"7e",x"50",x"c0"),
   960 => (x"49",x"bf",x"e8",x"f2"),
   961 => (x"bf",x"d8",x"ea",x"c2"),
   962 => (x"04",x"aa",x"71",x"4a"),
   963 => (x"cf",x"87",x"f4",x"fb"),
   964 => (x"f8",x"ff",x"ff",x"ff"),
   965 => (x"cc",x"f7",x"c2",x"4c"),
   966 => (x"c8",x"c0",x"05",x"bf"),
   967 => (x"e4",x"f2",x"c2",x"87"),
   968 => (x"fa",x"c1",x"02",x"bf"),
   969 => (x"d4",x"ea",x"c2",x"87"),
   970 => (x"f5",x"e6",x"49",x"bf"),
   971 => (x"d8",x"ea",x"c2",x"87"),
   972 => (x"48",x"a6",x"c4",x"58"),
   973 => (x"bf",x"d4",x"ea",x"c2"),
   974 => (x"e4",x"f2",x"c2",x"78"),
   975 => (x"db",x"c0",x"02",x"bf"),
   976 => (x"49",x"66",x"c4",x"87"),
   977 => (x"a9",x"74",x"99",x"74"),
   978 => (x"87",x"c8",x"c0",x"02"),
   979 => (x"c0",x"48",x"a6",x"c8"),
   980 => (x"87",x"e7",x"c0",x"78"),
   981 => (x"c1",x"48",x"a6",x"c8"),
   982 => (x"87",x"df",x"c0",x"78"),
   983 => (x"cf",x"49",x"66",x"c4"),
   984 => (x"a9",x"99",x"f8",x"ff"),
   985 => (x"87",x"c8",x"c0",x"02"),
   986 => (x"c0",x"48",x"a6",x"cc"),
   987 => (x"87",x"c5",x"c0",x"78"),
   988 => (x"c1",x"48",x"a6",x"cc"),
   989 => (x"48",x"a6",x"c8",x"78"),
   990 => (x"c8",x"78",x"66",x"cc"),
   991 => (x"de",x"c0",x"05",x"66"),
   992 => (x"49",x"66",x"c4",x"87"),
   993 => (x"f2",x"c2",x"89",x"c2"),
   994 => (x"c2",x"91",x"bf",x"dc"),
   995 => (x"48",x"bf",x"f8",x"f6"),
   996 => (x"ea",x"c2",x"80",x"71"),
   997 => (x"ea",x"c2",x"58",x"d4"),
   998 => (x"78",x"c0",x"48",x"d8"),
   999 => (x"c0",x"87",x"d4",x"f9"),
  1000 => (x"ff",x"ff",x"cf",x"48"),
  1001 => (x"f0",x"4c",x"f8",x"ff"),
  1002 => (x"26",x"4d",x"26",x"8e"),
  1003 => (x"26",x"4b",x"26",x"4c"),
  1004 => (x"00",x"00",x"00",x"4f"),
  1005 => (x"00",x"00",x"00",x"00"),
  1006 => (x"ff",x"ff",x"ff",x"ff"),
  1007 => (x"00",x"00",x"0f",x"c4"),
  1008 => (x"00",x"00",x"0f",x"d0"),
  1009 => (x"33",x"54",x"41",x"46"),
  1010 => (x"20",x"20",x"20",x"32"),
  1011 => (x"00",x"00",x"00",x"00"),
  1012 => (x"31",x"54",x"41",x"46"),
  1013 => (x"20",x"20",x"20",x"36"),
  1014 => (x"d4",x"ff",x"1e",x"00"),
  1015 => (x"78",x"ff",x"c3",x"48"),
  1016 => (x"4f",x"26",x"48",x"68"),
  1017 => (x"48",x"d4",x"ff",x"1e"),
  1018 => (x"ff",x"78",x"ff",x"c3"),
  1019 => (x"e1",x"c0",x"48",x"d0"),
  1020 => (x"48",x"d4",x"ff",x"78"),
  1021 => (x"4f",x"26",x"78",x"d4"),
  1022 => (x"48",x"d0",x"ff",x"1e"),
  1023 => (x"26",x"78",x"e0",x"c0"),
  1024 => (x"d4",x"ff",x"1e",x"4f"),
  1025 => (x"99",x"49",x"70",x"87"),
  1026 => (x"c0",x"87",x"c6",x"02"),
  1027 => (x"f1",x"05",x"a9",x"fb"),
  1028 => (x"26",x"48",x"71",x"87"),
  1029 => (x"5b",x"5e",x"0e",x"4f"),
  1030 => (x"4b",x"71",x"0e",x"5c"),
  1031 => (x"f8",x"fe",x"4c",x"c0"),
  1032 => (x"99",x"49",x"70",x"87"),
  1033 => (x"87",x"f9",x"c0",x"02"),
  1034 => (x"02",x"a9",x"ec",x"c0"),
  1035 => (x"c0",x"87",x"f2",x"c0"),
  1036 => (x"c0",x"02",x"a9",x"fb"),
  1037 => (x"66",x"cc",x"87",x"eb"),
  1038 => (x"c7",x"03",x"ac",x"b7"),
  1039 => (x"02",x"66",x"d0",x"87"),
  1040 => (x"53",x"71",x"87",x"c2"),
  1041 => (x"c2",x"02",x"99",x"71"),
  1042 => (x"fe",x"84",x"c1",x"87"),
  1043 => (x"49",x"70",x"87",x"cb"),
  1044 => (x"87",x"cd",x"02",x"99"),
  1045 => (x"02",x"a9",x"ec",x"c0"),
  1046 => (x"fb",x"c0",x"87",x"c7"),
  1047 => (x"d5",x"ff",x"05",x"a9"),
  1048 => (x"02",x"66",x"d0",x"87"),
  1049 => (x"97",x"c0",x"87",x"c3"),
  1050 => (x"a9",x"ec",x"c0",x"7b"),
  1051 => (x"74",x"87",x"c4",x"05"),
  1052 => (x"74",x"87",x"c5",x"4a"),
  1053 => (x"8a",x"0a",x"c0",x"4a"),
  1054 => (x"4c",x"26",x"48",x"72"),
  1055 => (x"4f",x"26",x"4b",x"26"),
  1056 => (x"87",x"d5",x"fd",x"1e"),
  1057 => (x"c0",x"4a",x"49",x"70"),
  1058 => (x"c9",x"04",x"aa",x"f0"),
  1059 => (x"aa",x"f9",x"c0",x"87"),
  1060 => (x"c0",x"87",x"c3",x"01"),
  1061 => (x"c1",x"c1",x"8a",x"f0"),
  1062 => (x"87",x"c9",x"04",x"aa"),
  1063 => (x"01",x"aa",x"da",x"c1"),
  1064 => (x"f7",x"c0",x"87",x"c3"),
  1065 => (x"26",x"48",x"72",x"8a"),
  1066 => (x"5b",x"5e",x"0e",x"4f"),
  1067 => (x"f8",x"0e",x"5d",x"5c"),
  1068 => (x"c0",x"4c",x"71",x"86"),
  1069 => (x"87",x"ec",x"fc",x"7e"),
  1070 => (x"c5",x"c1",x"4b",x"c0"),
  1071 => (x"49",x"bf",x"97",x"c8"),
  1072 => (x"cf",x"04",x"a9",x"c0"),
  1073 => (x"87",x"f9",x"fc",x"87"),
  1074 => (x"c5",x"c1",x"83",x"c1"),
  1075 => (x"49",x"bf",x"97",x"c8"),
  1076 => (x"87",x"f1",x"06",x"ab"),
  1077 => (x"97",x"c8",x"c5",x"c1"),
  1078 => (x"87",x"cf",x"02",x"bf"),
  1079 => (x"70",x"87",x"fa",x"fb"),
  1080 => (x"c6",x"02",x"99",x"49"),
  1081 => (x"a9",x"ec",x"c0",x"87"),
  1082 => (x"c0",x"87",x"f1",x"05"),
  1083 => (x"87",x"e9",x"fb",x"4b"),
  1084 => (x"e4",x"fb",x"4d",x"70"),
  1085 => (x"58",x"a6",x"c8",x"87"),
  1086 => (x"70",x"87",x"de",x"fb"),
  1087 => (x"c8",x"83",x"c1",x"4a"),
  1088 => (x"69",x"97",x"49",x"a4"),
  1089 => (x"da",x"05",x"ad",x"49"),
  1090 => (x"49",x"a4",x"c9",x"87"),
  1091 => (x"c4",x"49",x"69",x"97"),
  1092 => (x"ce",x"05",x"a9",x"66"),
  1093 => (x"49",x"a4",x"ca",x"87"),
  1094 => (x"aa",x"49",x"69",x"97"),
  1095 => (x"c1",x"87",x"c4",x"05"),
  1096 => (x"c0",x"87",x"d0",x"7e"),
  1097 => (x"c6",x"02",x"ad",x"ec"),
  1098 => (x"ad",x"fb",x"c0",x"87"),
  1099 => (x"c0",x"87",x"c4",x"05"),
  1100 => (x"6e",x"7e",x"c1",x"4b"),
  1101 => (x"87",x"f5",x"fe",x"02"),
  1102 => (x"73",x"87",x"fd",x"fa"),
  1103 => (x"26",x"8e",x"f8",x"48"),
  1104 => (x"26",x"4c",x"26",x"4d"),
  1105 => (x"00",x"4f",x"26",x"4b"),
  1106 => (x"1e",x"73",x"1e",x"00"),
  1107 => (x"c8",x"4b",x"d4",x"ff"),
  1108 => (x"d0",x"ff",x"4a",x"66"),
  1109 => (x"78",x"c5",x"c8",x"48"),
  1110 => (x"c1",x"48",x"d4",x"ff"),
  1111 => (x"7b",x"11",x"78",x"d4"),
  1112 => (x"f9",x"05",x"8a",x"c1"),
  1113 => (x"48",x"d0",x"ff",x"87"),
  1114 => (x"4b",x"26",x"78",x"c4"),
  1115 => (x"5e",x"0e",x"4f",x"26"),
  1116 => (x"0e",x"5d",x"5c",x"5b"),
  1117 => (x"7e",x"71",x"86",x"f8"),
  1118 => (x"f7",x"c2",x"1e",x"6e"),
  1119 => (x"df",x"ff",x"49",x"dc"),
  1120 => (x"86",x"c4",x"87",x"d7"),
  1121 => (x"c4",x"02",x"98",x"70"),
  1122 => (x"f4",x"c1",x"87",x"e4"),
  1123 => (x"6e",x"4c",x"bf",x"d0"),
  1124 => (x"87",x"d5",x"fc",x"49"),
  1125 => (x"70",x"58",x"a6",x"c8"),
  1126 => (x"87",x"c5",x"05",x"98"),
  1127 => (x"c1",x"48",x"a6",x"c4"),
  1128 => (x"48",x"d0",x"ff",x"78"),
  1129 => (x"d4",x"ff",x"78",x"c5"),
  1130 => (x"78",x"d5",x"c1",x"48"),
  1131 => (x"c1",x"49",x"66",x"c4"),
  1132 => (x"c1",x"31",x"c6",x"89"),
  1133 => (x"bf",x"97",x"c8",x"f4"),
  1134 => (x"b0",x"71",x"48",x"4a"),
  1135 => (x"78",x"08",x"d4",x"ff"),
  1136 => (x"c4",x"48",x"d0",x"ff"),
  1137 => (x"d8",x"f7",x"c2",x"78"),
  1138 => (x"d0",x"49",x"bf",x"97"),
  1139 => (x"87",x"dd",x"02",x"99"),
  1140 => (x"d4",x"ff",x"78",x"c5"),
  1141 => (x"78",x"d6",x"c1",x"48"),
  1142 => (x"d4",x"ff",x"4a",x"c0"),
  1143 => (x"78",x"ff",x"c3",x"48"),
  1144 => (x"e0",x"c0",x"82",x"c1"),
  1145 => (x"87",x"f2",x"04",x"aa"),
  1146 => (x"c4",x"48",x"d0",x"ff"),
  1147 => (x"48",x"d4",x"ff",x"78"),
  1148 => (x"ff",x"78",x"ff",x"c3"),
  1149 => (x"78",x"c5",x"48",x"d0"),
  1150 => (x"c1",x"48",x"d4",x"ff"),
  1151 => (x"78",x"c1",x"78",x"d3"),
  1152 => (x"c4",x"48",x"d0",x"ff"),
  1153 => (x"ac",x"b7",x"c0",x"78"),
  1154 => (x"87",x"cb",x"c2",x"06"),
  1155 => (x"bf",x"e4",x"f7",x"c2"),
  1156 => (x"7e",x"74",x"8c",x"4b"),
  1157 => (x"c1",x"02",x"9b",x"73"),
  1158 => (x"c0",x"c8",x"87",x"dd"),
  1159 => (x"b7",x"c0",x"8b",x"4d"),
  1160 => (x"87",x"c6",x"03",x"ab"),
  1161 => (x"4d",x"a3",x"c0",x"c8"),
  1162 => (x"f7",x"c2",x"4b",x"c0"),
  1163 => (x"49",x"bf",x"97",x"d8"),
  1164 => (x"cf",x"02",x"99",x"d0"),
  1165 => (x"c2",x"1e",x"c0",x"87"),
  1166 => (x"e2",x"49",x"dc",x"f7"),
  1167 => (x"86",x"c4",x"87",x"d9"),
  1168 => (x"87",x"d8",x"4c",x"70"),
  1169 => (x"1e",x"dc",x"ea",x"c2"),
  1170 => (x"49",x"dc",x"f7",x"c2"),
  1171 => (x"70",x"87",x"c8",x"e2"),
  1172 => (x"c2",x"1e",x"75",x"4c"),
  1173 => (x"fb",x"49",x"dc",x"ea"),
  1174 => (x"86",x"c8",x"87",x"ef"),
  1175 => (x"c5",x"05",x"9c",x"74"),
  1176 => (x"c1",x"48",x"c0",x"87"),
  1177 => (x"1e",x"c1",x"87",x"ca"),
  1178 => (x"49",x"dc",x"f7",x"c2"),
  1179 => (x"c4",x"87",x"cd",x"e0"),
  1180 => (x"05",x"9b",x"73",x"86"),
  1181 => (x"6e",x"87",x"e3",x"fe"),
  1182 => (x"ac",x"b7",x"c0",x"4c"),
  1183 => (x"c2",x"87",x"d1",x"06"),
  1184 => (x"c0",x"48",x"dc",x"f7"),
  1185 => (x"c0",x"80",x"d0",x"78"),
  1186 => (x"c2",x"80",x"f4",x"78"),
  1187 => (x"78",x"bf",x"e8",x"f7"),
  1188 => (x"01",x"ac",x"b7",x"c0"),
  1189 => (x"ff",x"87",x"f5",x"fd"),
  1190 => (x"78",x"c5",x"48",x"d0"),
  1191 => (x"c1",x"48",x"d4",x"ff"),
  1192 => (x"78",x"c0",x"78",x"d3"),
  1193 => (x"c4",x"48",x"d0",x"ff"),
  1194 => (x"c0",x"48",x"c1",x"78"),
  1195 => (x"48",x"c0",x"87",x"c2"),
  1196 => (x"4d",x"26",x"8e",x"f8"),
  1197 => (x"4b",x"26",x"4c",x"26"),
  1198 => (x"5e",x"0e",x"4f",x"26"),
  1199 => (x"0e",x"5d",x"5c",x"5b"),
  1200 => (x"4d",x"71",x"86",x"fc"),
  1201 => (x"ad",x"4c",x"4b",x"c0"),
  1202 => (x"87",x"e8",x"c0",x"04"),
  1203 => (x"1e",x"e9",x"c2",x"c1"),
  1204 => (x"c4",x"02",x"9c",x"74"),
  1205 => (x"c2",x"4a",x"c0",x"87"),
  1206 => (x"72",x"4a",x"c1",x"87"),
  1207 => (x"87",x"dd",x"eb",x"49"),
  1208 => (x"7e",x"70",x"86",x"c4"),
  1209 => (x"05",x"6e",x"83",x"c1"),
  1210 => (x"4b",x"75",x"87",x"c2"),
  1211 => (x"ab",x"75",x"84",x"c1"),
  1212 => (x"87",x"d8",x"ff",x"06"),
  1213 => (x"8e",x"fc",x"48",x"6e"),
  1214 => (x"4c",x"26",x"4d",x"26"),
  1215 => (x"4f",x"26",x"4b",x"26"),
  1216 => (x"5c",x"5b",x"5e",x"0e"),
  1217 => (x"cc",x"4b",x"71",x"0e"),
  1218 => (x"87",x"d8",x"02",x"66"),
  1219 => (x"8c",x"f0",x"c0",x"4c"),
  1220 => (x"74",x"87",x"d8",x"02"),
  1221 => (x"02",x"8a",x"c1",x"4a"),
  1222 => (x"02",x"8a",x"87",x"d1"),
  1223 => (x"02",x"8a",x"87",x"cd"),
  1224 => (x"87",x"d9",x"87",x"c9"),
  1225 => (x"c5",x"f9",x"49",x"73"),
  1226 => (x"74",x"87",x"d2",x"87"),
  1227 => (x"c1",x"49",x"c0",x"1e"),
  1228 => (x"74",x"87",x"fd",x"d9"),
  1229 => (x"c1",x"49",x"73",x"1e"),
  1230 => (x"c8",x"87",x"f5",x"d9"),
  1231 => (x"26",x"4c",x"26",x"86"),
  1232 => (x"0e",x"4f",x"26",x"4b"),
  1233 => (x"5d",x"5c",x"5b",x"5e"),
  1234 => (x"71",x"86",x"fc",x"0e"),
  1235 => (x"91",x"de",x"49",x"4c"),
  1236 => (x"4d",x"fc",x"f8",x"c2"),
  1237 => (x"6d",x"97",x"85",x"71"),
  1238 => (x"87",x"dc",x"c1",x"02"),
  1239 => (x"bf",x"ec",x"f8",x"c2"),
  1240 => (x"71",x"81",x"74",x"49"),
  1241 => (x"70",x"87",x"d3",x"fd"),
  1242 => (x"02",x"98",x"48",x"7e"),
  1243 => (x"c2",x"87",x"f2",x"c0"),
  1244 => (x"70",x"4b",x"f0",x"f8"),
  1245 => (x"fe",x"49",x"cb",x"4a"),
  1246 => (x"74",x"87",x"e9",x"f6"),
  1247 => (x"c1",x"93",x"cc",x"4b"),
  1248 => (x"c4",x"83",x"d4",x"f4"),
  1249 => (x"c4",x"cf",x"c1",x"83"),
  1250 => (x"c1",x"49",x"74",x"7b"),
  1251 => (x"75",x"87",x"e9",x"c4"),
  1252 => (x"cc",x"f4",x"c1",x"7b"),
  1253 => (x"1e",x"49",x"bf",x"97"),
  1254 => (x"49",x"f0",x"f8",x"c2"),
  1255 => (x"c4",x"87",x"e1",x"fd"),
  1256 => (x"c1",x"49",x"74",x"86"),
  1257 => (x"c0",x"87",x"d1",x"c4"),
  1258 => (x"ec",x"c5",x"c1",x"49"),
  1259 => (x"d4",x"f7",x"c2",x"87"),
  1260 => (x"49",x"50",x"c0",x"48"),
  1261 => (x"87",x"cb",x"e2",x"c0"),
  1262 => (x"4d",x"26",x"8e",x"fc"),
  1263 => (x"4b",x"26",x"4c",x"26"),
  1264 => (x"00",x"00",x"4f",x"26"),
  1265 => (x"64",x"61",x"6f",x"4c"),
  1266 => (x"2e",x"67",x"6e",x"69"),
  1267 => (x"1e",x"00",x"2e",x"2e"),
  1268 => (x"4b",x"71",x"1e",x"73"),
  1269 => (x"ec",x"f8",x"c2",x"49"),
  1270 => (x"fb",x"71",x"81",x"bf"),
  1271 => (x"4a",x"70",x"87",x"dc"),
  1272 => (x"87",x"c4",x"02",x"9a"),
  1273 => (x"87",x"db",x"e6",x"49"),
  1274 => (x"48",x"ec",x"f8",x"c2"),
  1275 => (x"49",x"73",x"78",x"c0"),
  1276 => (x"26",x"87",x"fa",x"c1"),
  1277 => (x"1e",x"4f",x"26",x"4b"),
  1278 => (x"4b",x"71",x"1e",x"73"),
  1279 => (x"02",x"4a",x"a3",x"c4"),
  1280 => (x"c1",x"87",x"d0",x"c1"),
  1281 => (x"87",x"dc",x"02",x"8a"),
  1282 => (x"f2",x"c0",x"02",x"8a"),
  1283 => (x"c1",x"05",x"8a",x"87"),
  1284 => (x"f8",x"c2",x"87",x"d3"),
  1285 => (x"c1",x"02",x"bf",x"ec"),
  1286 => (x"c1",x"48",x"87",x"cb"),
  1287 => (x"f0",x"f8",x"c2",x"88"),
  1288 => (x"87",x"c1",x"c1",x"58"),
  1289 => (x"bf",x"ec",x"f8",x"c2"),
  1290 => (x"c2",x"89",x"c6",x"49"),
  1291 => (x"c0",x"59",x"f0",x"f8"),
  1292 => (x"c0",x"03",x"a9",x"b7"),
  1293 => (x"f8",x"c2",x"87",x"ef"),
  1294 => (x"78",x"c0",x"48",x"ec"),
  1295 => (x"c2",x"87",x"e6",x"c0"),
  1296 => (x"02",x"bf",x"e8",x"f8"),
  1297 => (x"f8",x"c2",x"87",x"df"),
  1298 => (x"c1",x"48",x"bf",x"ec"),
  1299 => (x"f0",x"f8",x"c2",x"80"),
  1300 => (x"c2",x"87",x"d2",x"58"),
  1301 => (x"02",x"bf",x"e8",x"f8"),
  1302 => (x"f8",x"c2",x"87",x"cb"),
  1303 => (x"c6",x"48",x"bf",x"ec"),
  1304 => (x"f0",x"f8",x"c2",x"80"),
  1305 => (x"c4",x"49",x"73",x"58"),
  1306 => (x"26",x"4b",x"26",x"87"),
  1307 => (x"5b",x"5e",x"0e",x"4f"),
  1308 => (x"f0",x"0e",x"5d",x"5c"),
  1309 => (x"59",x"a6",x"d0",x"86"),
  1310 => (x"4d",x"dc",x"ea",x"c2"),
  1311 => (x"f8",x"c2",x"4c",x"c0"),
  1312 => (x"78",x"c1",x"48",x"e8"),
  1313 => (x"c0",x"48",x"a6",x"c8"),
  1314 => (x"c2",x"7e",x"75",x"78"),
  1315 => (x"48",x"bf",x"ec",x"f8"),
  1316 => (x"c1",x"06",x"a8",x"c0"),
  1317 => (x"a6",x"c8",x"87",x"c0"),
  1318 => (x"c2",x"7e",x"75",x"5c"),
  1319 => (x"98",x"48",x"dc",x"ea"),
  1320 => (x"87",x"f2",x"c0",x"02"),
  1321 => (x"c1",x"4d",x"66",x"c4"),
  1322 => (x"cc",x"1e",x"e9",x"c2"),
  1323 => (x"87",x"c4",x"02",x"66"),
  1324 => (x"87",x"c2",x"4c",x"c0"),
  1325 => (x"49",x"74",x"4c",x"c1"),
  1326 => (x"c4",x"87",x"c2",x"e4"),
  1327 => (x"c1",x"7e",x"70",x"86"),
  1328 => (x"48",x"66",x"c8",x"85"),
  1329 => (x"a6",x"cc",x"80",x"c1"),
  1330 => (x"ec",x"f8",x"c2",x"58"),
  1331 => (x"c5",x"03",x"ad",x"bf"),
  1332 => (x"ff",x"05",x"6e",x"87"),
  1333 => (x"4d",x"6e",x"87",x"d1"),
  1334 => (x"9d",x"75",x"4c",x"c0"),
  1335 => (x"87",x"dc",x"c3",x"02"),
  1336 => (x"1e",x"e9",x"c2",x"c1"),
  1337 => (x"c7",x"02",x"66",x"cc"),
  1338 => (x"48",x"a6",x"c8",x"87"),
  1339 => (x"87",x"c5",x"78",x"c0"),
  1340 => (x"c1",x"48",x"a6",x"c8"),
  1341 => (x"49",x"66",x"c8",x"78"),
  1342 => (x"c4",x"87",x"c2",x"e3"),
  1343 => (x"48",x"7e",x"70",x"86"),
  1344 => (x"e4",x"c2",x"02",x"98"),
  1345 => (x"81",x"cb",x"49",x"87"),
  1346 => (x"d0",x"49",x"69",x"97"),
  1347 => (x"d4",x"c1",x"02",x"99"),
  1348 => (x"cc",x"49",x"74",x"87"),
  1349 => (x"d4",x"f4",x"c1",x"91"),
  1350 => (x"cf",x"cf",x"c1",x"81"),
  1351 => (x"c3",x"81",x"c8",x"79"),
  1352 => (x"49",x"74",x"51",x"ff"),
  1353 => (x"f8",x"c2",x"91",x"de"),
  1354 => (x"85",x"71",x"4d",x"fc"),
  1355 => (x"7d",x"97",x"c1",x"c2"),
  1356 => (x"c0",x"49",x"a5",x"c1"),
  1357 => (x"f2",x"c2",x"51",x"e0"),
  1358 => (x"02",x"bf",x"97",x"ec"),
  1359 => (x"84",x"c1",x"87",x"d2"),
  1360 => (x"c2",x"4b",x"a5",x"c2"),
  1361 => (x"db",x"4a",x"ec",x"f2"),
  1362 => (x"d7",x"ef",x"fe",x"49"),
  1363 => (x"87",x"d9",x"c1",x"87"),
  1364 => (x"c0",x"49",x"a5",x"cd"),
  1365 => (x"c2",x"84",x"c1",x"51"),
  1366 => (x"4a",x"6e",x"4b",x"a5"),
  1367 => (x"ef",x"fe",x"49",x"cb"),
  1368 => (x"c4",x"c1",x"87",x"c2"),
  1369 => (x"cc",x"49",x"74",x"87"),
  1370 => (x"d4",x"f4",x"c1",x"91"),
  1371 => (x"c3",x"cd",x"c1",x"81"),
  1372 => (x"ec",x"f2",x"c2",x"79"),
  1373 => (x"d8",x"02",x"bf",x"97"),
  1374 => (x"de",x"49",x"74",x"87"),
  1375 => (x"c2",x"84",x"c1",x"91"),
  1376 => (x"71",x"4b",x"fc",x"f8"),
  1377 => (x"ec",x"f2",x"c2",x"83"),
  1378 => (x"fe",x"49",x"dd",x"4a"),
  1379 => (x"d8",x"87",x"d5",x"ee"),
  1380 => (x"de",x"4b",x"74",x"87"),
  1381 => (x"fc",x"f8",x"c2",x"93"),
  1382 => (x"49",x"a3",x"cb",x"83"),
  1383 => (x"84",x"c1",x"51",x"c0"),
  1384 => (x"cb",x"4a",x"6e",x"73"),
  1385 => (x"fb",x"ed",x"fe",x"49"),
  1386 => (x"48",x"66",x"c8",x"87"),
  1387 => (x"a6",x"cc",x"80",x"c1"),
  1388 => (x"03",x"ac",x"c7",x"58"),
  1389 => (x"6e",x"87",x"c5",x"c0"),
  1390 => (x"87",x"e4",x"fc",x"05"),
  1391 => (x"c0",x"03",x"ac",x"c7"),
  1392 => (x"f8",x"c2",x"87",x"e4"),
  1393 => (x"78",x"c0",x"48",x"e8"),
  1394 => (x"91",x"cc",x"49",x"74"),
  1395 => (x"81",x"d4",x"f4",x"c1"),
  1396 => (x"79",x"c3",x"cd",x"c1"),
  1397 => (x"91",x"de",x"49",x"74"),
  1398 => (x"81",x"fc",x"f8",x"c2"),
  1399 => (x"84",x"c1",x"51",x"c0"),
  1400 => (x"ff",x"04",x"ac",x"c7"),
  1401 => (x"f5",x"c1",x"87",x"dc"),
  1402 => (x"50",x"c0",x"48",x"f0"),
  1403 => (x"d9",x"c1",x"80",x"f7"),
  1404 => (x"d8",x"c1",x"40",x"dd"),
  1405 => (x"80",x"c8",x"78",x"d0"),
  1406 => (x"78",x"f7",x"cf",x"c1"),
  1407 => (x"c0",x"49",x"66",x"cc"),
  1408 => (x"f0",x"87",x"f5",x"fa"),
  1409 => (x"26",x"4d",x"26",x"8e"),
  1410 => (x"26",x"4b",x"26",x"4c"),
  1411 => (x"00",x"00",x"00",x"4f"),
  1412 => (x"61",x"42",x"20",x"80"),
  1413 => (x"1e",x"00",x"6b",x"63"),
  1414 => (x"4b",x"71",x"1e",x"73"),
  1415 => (x"c1",x"91",x"cc",x"49"),
  1416 => (x"c8",x"81",x"d4",x"f4"),
  1417 => (x"f4",x"c1",x"4a",x"a1"),
  1418 => (x"50",x"12",x"48",x"c8"),
  1419 => (x"c1",x"4a",x"a1",x"c9"),
  1420 => (x"12",x"48",x"c8",x"c5"),
  1421 => (x"c1",x"81",x"ca",x"50"),
  1422 => (x"11",x"48",x"cc",x"f4"),
  1423 => (x"cc",x"f4",x"c1",x"50"),
  1424 => (x"1e",x"49",x"bf",x"97"),
  1425 => (x"f7",x"f2",x"49",x"c0"),
  1426 => (x"f8",x"49",x"73",x"87"),
  1427 => (x"8e",x"fc",x"87",x"df"),
  1428 => (x"4f",x"26",x"4b",x"26"),
  1429 => (x"c0",x"49",x"c0",x"1e"),
  1430 => (x"26",x"87",x"fe",x"fa"),
  1431 => (x"4a",x"71",x"1e",x"4f"),
  1432 => (x"c1",x"91",x"cc",x"49"),
  1433 => (x"c8",x"81",x"d4",x"f4"),
  1434 => (x"d4",x"f7",x"c2",x"81"),
  1435 => (x"c0",x"50",x"11",x"48"),
  1436 => (x"fe",x"49",x"a2",x"f0"),
  1437 => (x"c0",x"87",x"d5",x"e8"),
  1438 => (x"87",x"c7",x"d7",x"49"),
  1439 => (x"ff",x"1e",x"4f",x"26"),
  1440 => (x"ff",x"c3",x"4a",x"d4"),
  1441 => (x"48",x"d0",x"ff",x"7a"),
  1442 => (x"de",x"78",x"e1",x"c0"),
  1443 => (x"48",x"7a",x"71",x"7a"),
  1444 => (x"70",x"28",x"b7",x"c8"),
  1445 => (x"d0",x"48",x"71",x"7a"),
  1446 => (x"7a",x"70",x"28",x"b7"),
  1447 => (x"b7",x"d8",x"48",x"71"),
  1448 => (x"ff",x"7a",x"70",x"28"),
  1449 => (x"e0",x"c0",x"48",x"d0"),
  1450 => (x"0e",x"4f",x"26",x"78"),
  1451 => (x"5d",x"5c",x"5b",x"5e"),
  1452 => (x"71",x"86",x"f4",x"0e"),
  1453 => (x"91",x"cc",x"49",x"4d"),
  1454 => (x"81",x"d4",x"f4",x"c1"),
  1455 => (x"ca",x"4a",x"a1",x"c8"),
  1456 => (x"a6",x"c4",x"7e",x"a1"),
  1457 => (x"d0",x"f7",x"c2",x"48"),
  1458 => (x"97",x"6e",x"78",x"bf"),
  1459 => (x"66",x"c4",x"4b",x"bf"),
  1460 => (x"12",x"2c",x"73",x"4c"),
  1461 => (x"58",x"a6",x"cc",x"48"),
  1462 => (x"84",x"c1",x"9c",x"70"),
  1463 => (x"69",x"97",x"81",x"c9"),
  1464 => (x"04",x"ac",x"b7",x"49"),
  1465 => (x"4c",x"c0",x"87",x"c2"),
  1466 => (x"4a",x"bf",x"97",x"6e"),
  1467 => (x"72",x"49",x"66",x"c8"),
  1468 => (x"c4",x"b9",x"ff",x"31"),
  1469 => (x"48",x"74",x"99",x"66"),
  1470 => (x"4a",x"70",x"30",x"72"),
  1471 => (x"d4",x"f7",x"c2",x"b1"),
  1472 => (x"f9",x"fd",x"71",x"59"),
  1473 => (x"c2",x"1e",x"c7",x"87"),
  1474 => (x"1e",x"bf",x"e4",x"f8"),
  1475 => (x"1e",x"d4",x"f4",x"c1"),
  1476 => (x"97",x"d4",x"f7",x"c2"),
  1477 => (x"f4",x"c1",x"49",x"bf"),
  1478 => (x"c0",x"49",x"75",x"87"),
  1479 => (x"e8",x"87",x"d9",x"f6"),
  1480 => (x"26",x"4d",x"26",x"8e"),
  1481 => (x"26",x"4b",x"26",x"4c"),
  1482 => (x"1e",x"73",x"1e",x"4f"),
  1483 => (x"fd",x"49",x"4b",x"71"),
  1484 => (x"49",x"73",x"87",x"f9"),
  1485 => (x"26",x"87",x"f4",x"fd"),
  1486 => (x"1e",x"4f",x"26",x"4b"),
  1487 => (x"4b",x"71",x"1e",x"73"),
  1488 => (x"02",x"4a",x"a3",x"c2"),
  1489 => (x"8a",x"c1",x"87",x"d6"),
  1490 => (x"87",x"e2",x"c0",x"05"),
  1491 => (x"bf",x"e4",x"f8",x"c2"),
  1492 => (x"48",x"87",x"db",x"02"),
  1493 => (x"f8",x"c2",x"88",x"c1"),
  1494 => (x"87",x"d2",x"58",x"e8"),
  1495 => (x"bf",x"e8",x"f8",x"c2"),
  1496 => (x"c2",x"87",x"cb",x"02"),
  1497 => (x"48",x"bf",x"e4",x"f8"),
  1498 => (x"f8",x"c2",x"80",x"c1"),
  1499 => (x"1e",x"c7",x"58",x"e8"),
  1500 => (x"bf",x"e4",x"f8",x"c2"),
  1501 => (x"d4",x"f4",x"c1",x"1e"),
  1502 => (x"d4",x"f7",x"c2",x"1e"),
  1503 => (x"cc",x"49",x"bf",x"97"),
  1504 => (x"c0",x"49",x"73",x"87"),
  1505 => (x"f4",x"87",x"f1",x"f4"),
  1506 => (x"26",x"4b",x"26",x"8e"),
  1507 => (x"5b",x"5e",x"0e",x"4f"),
  1508 => (x"ff",x"0e",x"5d",x"5c"),
  1509 => (x"e4",x"c0",x"86",x"cc"),
  1510 => (x"a6",x"cc",x"59",x"a6"),
  1511 => (x"c4",x"78",x"c0",x"48"),
  1512 => (x"c4",x"78",x"c0",x"80"),
  1513 => (x"66",x"c8",x"c1",x"80"),
  1514 => (x"c1",x"80",x"c4",x"78"),
  1515 => (x"c1",x"80",x"c4",x"78"),
  1516 => (x"e8",x"f8",x"c2",x"78"),
  1517 => (x"e0",x"78",x"c1",x"48"),
  1518 => (x"c4",x"e1",x"87",x"ea"),
  1519 => (x"87",x"d9",x"e0",x"87"),
  1520 => (x"fb",x"c0",x"4c",x"70"),
  1521 => (x"f3",x"c1",x"02",x"ac"),
  1522 => (x"66",x"e0",x"c0",x"87"),
  1523 => (x"87",x"e8",x"c1",x"05"),
  1524 => (x"4a",x"66",x"c4",x"c1"),
  1525 => (x"7e",x"6a",x"82",x"c4"),
  1526 => (x"48",x"e4",x"f0",x"c1"),
  1527 => (x"41",x"20",x"49",x"6e"),
  1528 => (x"51",x"10",x"41",x"20"),
  1529 => (x"48",x"66",x"c4",x"c1"),
  1530 => (x"78",x"d7",x"d8",x"c1"),
  1531 => (x"81",x"c7",x"49",x"6a"),
  1532 => (x"c4",x"c1",x"51",x"74"),
  1533 => (x"81",x"c8",x"49",x"66"),
  1534 => (x"a6",x"d8",x"51",x"c1"),
  1535 => (x"c1",x"78",x"c2",x"48"),
  1536 => (x"c9",x"49",x"66",x"c4"),
  1537 => (x"c1",x"51",x"c0",x"81"),
  1538 => (x"ca",x"49",x"66",x"c4"),
  1539 => (x"c1",x"51",x"c0",x"81"),
  1540 => (x"6a",x"1e",x"d8",x"1e"),
  1541 => (x"ff",x"81",x"c8",x"49"),
  1542 => (x"c8",x"87",x"fa",x"df"),
  1543 => (x"66",x"c8",x"c1",x"86"),
  1544 => (x"01",x"a8",x"c0",x"48"),
  1545 => (x"a6",x"d0",x"87",x"c7"),
  1546 => (x"cf",x"78",x"c1",x"48"),
  1547 => (x"66",x"c8",x"c1",x"87"),
  1548 => (x"d8",x"88",x"c1",x"48"),
  1549 => (x"87",x"c4",x"58",x"a6"),
  1550 => (x"87",x"c5",x"df",x"ff"),
  1551 => (x"cd",x"02",x"9c",x"74"),
  1552 => (x"66",x"d0",x"87",x"da"),
  1553 => (x"66",x"cc",x"c1",x"48"),
  1554 => (x"cf",x"cd",x"03",x"a8"),
  1555 => (x"48",x"a6",x"c8",x"87"),
  1556 => (x"ff",x"7e",x"78",x"c0"),
  1557 => (x"70",x"87",x"c2",x"de"),
  1558 => (x"ac",x"d0",x"c1",x"4c"),
  1559 => (x"87",x"e7",x"c2",x"05"),
  1560 => (x"6e",x"48",x"a6",x"c4"),
  1561 => (x"87",x"d8",x"e0",x"78"),
  1562 => (x"cc",x"48",x"7e",x"70"),
  1563 => (x"c5",x"06",x"a8",x"66"),
  1564 => (x"48",x"a6",x"cc",x"87"),
  1565 => (x"dd",x"ff",x"78",x"6e"),
  1566 => (x"4c",x"70",x"87",x"df"),
  1567 => (x"05",x"ac",x"ec",x"c0"),
  1568 => (x"d0",x"87",x"ee",x"c1"),
  1569 => (x"91",x"cc",x"49",x"66"),
  1570 => (x"81",x"66",x"c4",x"c1"),
  1571 => (x"6a",x"4a",x"a1",x"c4"),
  1572 => (x"4a",x"a1",x"c8",x"4d"),
  1573 => (x"d9",x"c1",x"52",x"6e"),
  1574 => (x"dc",x"ff",x"79",x"dd"),
  1575 => (x"4c",x"70",x"87",x"fb"),
  1576 => (x"87",x"d9",x"02",x"9c"),
  1577 => (x"02",x"ac",x"fb",x"c0"),
  1578 => (x"55",x"74",x"87",x"d3"),
  1579 => (x"87",x"e9",x"dc",x"ff"),
  1580 => (x"02",x"9c",x"4c",x"70"),
  1581 => (x"fb",x"c0",x"87",x"c7"),
  1582 => (x"ed",x"ff",x"05",x"ac"),
  1583 => (x"55",x"e0",x"c0",x"87"),
  1584 => (x"c0",x"55",x"c1",x"c2"),
  1585 => (x"e0",x"c0",x"7d",x"97"),
  1586 => (x"66",x"c4",x"48",x"66"),
  1587 => (x"87",x"db",x"05",x"a8"),
  1588 => (x"d4",x"48",x"66",x"d0"),
  1589 => (x"ca",x"04",x"a8",x"66"),
  1590 => (x"48",x"66",x"d0",x"87"),
  1591 => (x"a6",x"d4",x"80",x"c1"),
  1592 => (x"d4",x"87",x"c8",x"58"),
  1593 => (x"88",x"c1",x"48",x"66"),
  1594 => (x"ff",x"58",x"a6",x"d8"),
  1595 => (x"70",x"87",x"ea",x"db"),
  1596 => (x"ac",x"d0",x"c1",x"4c"),
  1597 => (x"dc",x"87",x"c9",x"05"),
  1598 => (x"80",x"c1",x"48",x"66"),
  1599 => (x"58",x"a6",x"e0",x"c0"),
  1600 => (x"02",x"ac",x"d0",x"c1"),
  1601 => (x"6e",x"87",x"d9",x"fd"),
  1602 => (x"66",x"e0",x"c0",x"48"),
  1603 => (x"eb",x"c9",x"05",x"a8"),
  1604 => (x"a6",x"e4",x"c0",x"87"),
  1605 => (x"74",x"78",x"c0",x"48"),
  1606 => (x"88",x"fb",x"c0",x"48"),
  1607 => (x"70",x"58",x"a6",x"c8"),
  1608 => (x"dd",x"c9",x"02",x"98"),
  1609 => (x"88",x"cb",x"48",x"87"),
  1610 => (x"70",x"58",x"a6",x"c8"),
  1611 => (x"cf",x"c1",x"02",x"98"),
  1612 => (x"88",x"c9",x"48",x"87"),
  1613 => (x"70",x"58",x"a6",x"c8"),
  1614 => (x"ff",x"c3",x"02",x"98"),
  1615 => (x"88",x"c4",x"48",x"87"),
  1616 => (x"70",x"58",x"a6",x"c8"),
  1617 => (x"87",x"cf",x"02",x"98"),
  1618 => (x"c8",x"88",x"c1",x"48"),
  1619 => (x"98",x"70",x"58",x"a6"),
  1620 => (x"87",x"e8",x"c3",x"02"),
  1621 => (x"c8",x"87",x"dc",x"c8"),
  1622 => (x"f0",x"c0",x"48",x"a6"),
  1623 => (x"f8",x"d9",x"ff",x"78"),
  1624 => (x"c0",x"4c",x"70",x"87"),
  1625 => (x"c0",x"02",x"ac",x"ec"),
  1626 => (x"a6",x"cc",x"87",x"c3"),
  1627 => (x"ac",x"ec",x"c0",x"5c"),
  1628 => (x"ff",x"87",x"cd",x"02"),
  1629 => (x"70",x"87",x"e2",x"d9"),
  1630 => (x"ac",x"ec",x"c0",x"4c"),
  1631 => (x"87",x"f3",x"ff",x"05"),
  1632 => (x"02",x"ac",x"ec",x"c0"),
  1633 => (x"ff",x"87",x"c4",x"c0"),
  1634 => (x"c0",x"87",x"ce",x"d9"),
  1635 => (x"d8",x"1e",x"ca",x"1e"),
  1636 => (x"91",x"cc",x"49",x"66"),
  1637 => (x"48",x"66",x"cc",x"c1"),
  1638 => (x"a6",x"cc",x"80",x"71"),
  1639 => (x"48",x"66",x"c8",x"58"),
  1640 => (x"a6",x"d0",x"80",x"c4"),
  1641 => (x"bf",x"66",x"cc",x"58"),
  1642 => (x"e8",x"d9",x"ff",x"49"),
  1643 => (x"de",x"1e",x"c1",x"87"),
  1644 => (x"bf",x"66",x"d4",x"1e"),
  1645 => (x"dc",x"d9",x"ff",x"49"),
  1646 => (x"70",x"86",x"d0",x"87"),
  1647 => (x"08",x"c0",x"48",x"49"),
  1648 => (x"a6",x"ec",x"c0",x"88"),
  1649 => (x"06",x"a8",x"c0",x"58"),
  1650 => (x"c0",x"87",x"ee",x"c0"),
  1651 => (x"dd",x"48",x"66",x"e8"),
  1652 => (x"e4",x"c0",x"03",x"a8"),
  1653 => (x"bf",x"66",x"c4",x"87"),
  1654 => (x"66",x"e8",x"c0",x"49"),
  1655 => (x"51",x"e0",x"c0",x"81"),
  1656 => (x"49",x"66",x"e8",x"c0"),
  1657 => (x"66",x"c4",x"81",x"c1"),
  1658 => (x"c1",x"c2",x"81",x"bf"),
  1659 => (x"66",x"e8",x"c0",x"51"),
  1660 => (x"c4",x"81",x"c2",x"49"),
  1661 => (x"c0",x"81",x"bf",x"66"),
  1662 => (x"c1",x"48",x"6e",x"51"),
  1663 => (x"6e",x"78",x"d7",x"d8"),
  1664 => (x"d8",x"81",x"c8",x"49"),
  1665 => (x"49",x"6e",x"51",x"66"),
  1666 => (x"66",x"dc",x"81",x"c9"),
  1667 => (x"ca",x"49",x"6e",x"51"),
  1668 => (x"51",x"66",x"c8",x"81"),
  1669 => (x"c1",x"48",x"66",x"d8"),
  1670 => (x"58",x"a6",x"dc",x"80"),
  1671 => (x"d4",x"48",x"66",x"d0"),
  1672 => (x"c0",x"04",x"a8",x"66"),
  1673 => (x"66",x"d0",x"87",x"cb"),
  1674 => (x"d4",x"80",x"c1",x"48"),
  1675 => (x"d1",x"c5",x"58",x"a6"),
  1676 => (x"48",x"66",x"d4",x"87"),
  1677 => (x"a6",x"d8",x"88",x"c1"),
  1678 => (x"87",x"c6",x"c5",x"58"),
  1679 => (x"87",x"c0",x"d9",x"ff"),
  1680 => (x"58",x"a6",x"ec",x"c0"),
  1681 => (x"87",x"f8",x"d8",x"ff"),
  1682 => (x"58",x"a6",x"f0",x"c0"),
  1683 => (x"05",x"a8",x"ec",x"c0"),
  1684 => (x"a6",x"87",x"c9",x"c0"),
  1685 => (x"66",x"e8",x"c0",x"48"),
  1686 => (x"87",x"c4",x"c0",x"78"),
  1687 => (x"87",x"f9",x"d5",x"ff"),
  1688 => (x"cc",x"49",x"66",x"d0"),
  1689 => (x"66",x"c4",x"c1",x"91"),
  1690 => (x"c8",x"80",x"71",x"48"),
  1691 => (x"66",x"c4",x"58",x"a6"),
  1692 => (x"c4",x"82",x"c8",x"4a"),
  1693 => (x"81",x"ca",x"49",x"66"),
  1694 => (x"51",x"66",x"e8",x"c0"),
  1695 => (x"49",x"66",x"ec",x"c0"),
  1696 => (x"e8",x"c0",x"81",x"c1"),
  1697 => (x"48",x"c1",x"89",x"66"),
  1698 => (x"49",x"70",x"30",x"71"),
  1699 => (x"97",x"71",x"89",x"c1"),
  1700 => (x"d0",x"f7",x"c2",x"7a"),
  1701 => (x"e8",x"c0",x"49",x"bf"),
  1702 => (x"6a",x"97",x"29",x"66"),
  1703 => (x"98",x"71",x"48",x"4a"),
  1704 => (x"58",x"a6",x"f4",x"c0"),
  1705 => (x"c4",x"48",x"66",x"c4"),
  1706 => (x"58",x"a6",x"cc",x"80"),
  1707 => (x"4d",x"bf",x"66",x"c8"),
  1708 => (x"48",x"66",x"e0",x"c0"),
  1709 => (x"c0",x"02",x"a8",x"6e"),
  1710 => (x"7e",x"c0",x"87",x"c5"),
  1711 => (x"c1",x"87",x"c2",x"c0"),
  1712 => (x"c0",x"1e",x"6e",x"7e"),
  1713 => (x"49",x"75",x"1e",x"e0"),
  1714 => (x"87",x"c9",x"d5",x"ff"),
  1715 => (x"4c",x"70",x"86",x"c8"),
  1716 => (x"06",x"ac",x"b7",x"c0"),
  1717 => (x"74",x"87",x"d4",x"c1"),
  1718 => (x"bf",x"66",x"c8",x"85"),
  1719 => (x"81",x"e0",x"c0",x"49"),
  1720 => (x"c1",x"4b",x"89",x"75"),
  1721 => (x"71",x"4a",x"f0",x"f0"),
  1722 => (x"87",x"f8",x"d8",x"fe"),
  1723 => (x"7e",x"75",x"85",x"c2"),
  1724 => (x"48",x"66",x"e4",x"c0"),
  1725 => (x"e8",x"c0",x"80",x"c1"),
  1726 => (x"f0",x"c0",x"58",x"a6"),
  1727 => (x"81",x"c1",x"49",x"66"),
  1728 => (x"c0",x"02",x"a9",x"70"),
  1729 => (x"4d",x"c0",x"87",x"c5"),
  1730 => (x"c1",x"87",x"c2",x"c0"),
  1731 => (x"cc",x"1e",x"75",x"4d"),
  1732 => (x"c0",x"49",x"bf",x"66"),
  1733 => (x"66",x"c4",x"81",x"e0"),
  1734 => (x"c8",x"1e",x"71",x"89"),
  1735 => (x"d3",x"ff",x"49",x"66"),
  1736 => (x"86",x"c8",x"87",x"f3"),
  1737 => (x"01",x"a8",x"b7",x"c0"),
  1738 => (x"c0",x"87",x"c5",x"ff"),
  1739 => (x"c0",x"02",x"66",x"e4"),
  1740 => (x"66",x"c4",x"87",x"d3"),
  1741 => (x"c0",x"81",x"c9",x"49"),
  1742 => (x"c4",x"51",x"66",x"e4"),
  1743 => (x"da",x"c1",x"48",x"66"),
  1744 => (x"ce",x"c0",x"78",x"eb"),
  1745 => (x"49",x"66",x"c4",x"87"),
  1746 => (x"51",x"c2",x"81",x"c9"),
  1747 => (x"c1",x"48",x"66",x"c4"),
  1748 => (x"d0",x"78",x"e9",x"dc"),
  1749 => (x"66",x"d4",x"48",x"66"),
  1750 => (x"cb",x"c0",x"04",x"a8"),
  1751 => (x"48",x"66",x"d0",x"87"),
  1752 => (x"a6",x"d4",x"80",x"c1"),
  1753 => (x"87",x"da",x"c0",x"58"),
  1754 => (x"c1",x"48",x"66",x"d4"),
  1755 => (x"58",x"a6",x"d8",x"88"),
  1756 => (x"ff",x"87",x"cf",x"c0"),
  1757 => (x"70",x"87",x"ca",x"d2"),
  1758 => (x"87",x"c6",x"c0",x"4c"),
  1759 => (x"87",x"c1",x"d2",x"ff"),
  1760 => (x"66",x"dc",x"4c",x"70"),
  1761 => (x"c0",x"80",x"c1",x"48"),
  1762 => (x"74",x"58",x"a6",x"e0"),
  1763 => (x"cb",x"c0",x"02",x"9c"),
  1764 => (x"48",x"66",x"d0",x"87"),
  1765 => (x"a8",x"66",x"cc",x"c1"),
  1766 => (x"87",x"f1",x"f2",x"04"),
  1767 => (x"c7",x"48",x"66",x"d0"),
  1768 => (x"e1",x"c0",x"03",x"a8"),
  1769 => (x"4c",x"66",x"d0",x"87"),
  1770 => (x"48",x"e8",x"f8",x"c2"),
  1771 => (x"49",x"74",x"78",x"c0"),
  1772 => (x"c4",x"c1",x"91",x"cc"),
  1773 => (x"a1",x"c4",x"81",x"66"),
  1774 => (x"c0",x"4a",x"6a",x"4a"),
  1775 => (x"84",x"c1",x"79",x"52"),
  1776 => (x"ff",x"04",x"ac",x"c7"),
  1777 => (x"e0",x"c0",x"87",x"e2"),
  1778 => (x"e2",x"c0",x"02",x"66"),
  1779 => (x"66",x"c4",x"c1",x"87"),
  1780 => (x"81",x"d4",x"c1",x"49"),
  1781 => (x"4a",x"66",x"c4",x"c1"),
  1782 => (x"c0",x"82",x"dc",x"c1"),
  1783 => (x"dd",x"d9",x"c1",x"52"),
  1784 => (x"66",x"c4",x"c1",x"79"),
  1785 => (x"81",x"d8",x"c1",x"49"),
  1786 => (x"79",x"f4",x"f0",x"c1"),
  1787 => (x"c1",x"87",x"d6",x"c0"),
  1788 => (x"c1",x"49",x"66",x"c4"),
  1789 => (x"c4",x"c1",x"81",x"d4"),
  1790 => (x"d8",x"c1",x"4a",x"66"),
  1791 => (x"fc",x"f0",x"c1",x"82"),
  1792 => (x"d4",x"d9",x"c1",x"7a"),
  1793 => (x"66",x"c4",x"c1",x"79"),
  1794 => (x"81",x"e0",x"c1",x"49"),
  1795 => (x"79",x"fb",x"dc",x"c1"),
  1796 => (x"87",x"e4",x"cf",x"ff"),
  1797 => (x"ff",x"48",x"66",x"cc"),
  1798 => (x"4d",x"26",x"8e",x"cc"),
  1799 => (x"4b",x"26",x"4c",x"26"),
  1800 => (x"00",x"00",x"4f",x"26"),
  1801 => (x"64",x"61",x"6f",x"4c"),
  1802 => (x"20",x"2e",x"2a",x"20"),
  1803 => (x"00",x"00",x"00",x"00"),
  1804 => (x"00",x"00",x"20",x"3a"),
  1805 => (x"61",x"42",x"20",x"80"),
  1806 => (x"00",x"00",x"6b",x"63"),
  1807 => (x"78",x"45",x"20",x"80"),
  1808 => (x"1e",x"00",x"74",x"69"),
  1809 => (x"f8",x"c2",x"1e",x"c7"),
  1810 => (x"c1",x"1e",x"bf",x"e4"),
  1811 => (x"c2",x"1e",x"d4",x"f4"),
  1812 => (x"bf",x"97",x"d4",x"f7"),
  1813 => (x"87",x"f5",x"ec",x"49"),
  1814 => (x"49",x"d4",x"f4",x"c1"),
  1815 => (x"87",x"e6",x"e2",x"c0"),
  1816 => (x"4f",x"26",x"8e",x"f4"),
  1817 => (x"c8",x"1e",x"73",x"1e"),
  1818 => (x"f5",x"c1",x"87",x"c3"),
  1819 => (x"f3",x"c1",x"48",x"ec"),
  1820 => (x"e8",x"fe",x"78",x"f4"),
  1821 => (x"e2",x"c0",x"49",x"a0"),
  1822 => (x"49",x"c7",x"87",x"cc"),
  1823 => (x"87",x"f8",x"e0",x"c0"),
  1824 => (x"e2",x"c0",x"49",x"c1"),
  1825 => (x"d4",x"ff",x"87",x"d3"),
  1826 => (x"78",x"ff",x"c3",x"48"),
  1827 => (x"48",x"f0",x"f8",x"c2"),
  1828 => (x"dd",x"fe",x"50",x"c0"),
  1829 => (x"98",x"70",x"87",x"da"),
  1830 => (x"fe",x"87",x"cd",x"02"),
  1831 => (x"70",x"87",x"d6",x"e7"),
  1832 => (x"87",x"c4",x"02",x"98"),
  1833 => (x"87",x"c2",x"4a",x"c1"),
  1834 => (x"9a",x"72",x"4a",x"c0"),
  1835 => (x"c1",x"87",x"c8",x"02"),
  1836 => (x"fe",x"49",x"c0",x"f4"),
  1837 => (x"c2",x"87",x"f0",x"cf"),
  1838 => (x"c0",x"48",x"e4",x"f8"),
  1839 => (x"d4",x"f7",x"c2",x"78"),
  1840 => (x"49",x"50",x"c0",x"48"),
  1841 => (x"c0",x"87",x"fc",x"fd"),
  1842 => (x"70",x"87",x"ea",x"f5"),
  1843 => (x"cb",x"02",x"9b",x"4b"),
  1844 => (x"f0",x"f5",x"c1",x"87"),
  1845 => (x"df",x"49",x"c7",x"5b"),
  1846 => (x"87",x"c6",x"87",x"de"),
  1847 => (x"e0",x"c0",x"49",x"c0"),
  1848 => (x"c2",x"c3",x"87",x"f7"),
  1849 => (x"d8",x"e2",x"c0",x"87"),
  1850 => (x"ec",x"ef",x"c0",x"87"),
  1851 => (x"87",x"f5",x"ff",x"87"),
  1852 => (x"4f",x"26",x"4b",x"26"),
  1853 => (x"74",x"6f",x"6f",x"42"),
  1854 => (x"2e",x"67",x"6e",x"69"),
  1855 => (x"00",x"00",x"2e",x"2e"),
  1856 => (x"4f",x"20",x"44",x"53"),
  1857 => (x"00",x"00",x"00",x"4b"),
  1858 => (x"00",x"00",x"00",x"00"),
  1859 => (x"00",x"00",x"00",x"00"),
  1860 => (x"00",x"00",x"00",x"01"),
  1861 => (x"00",x"00",x"13",x"43"),
  1862 => (x"00",x"00",x"2e",x"3c"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"13",x"43"),
  1865 => (x"00",x"00",x"2e",x"5a"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"00",x"00",x"13",x"43"),
  1868 => (x"00",x"00",x"2e",x"78"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"13",x"43"),
  1871 => (x"00",x"00",x"2e",x"96"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"13",x"43"),
  1874 => (x"00",x"00",x"2e",x"b4"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"13",x"43"),
  1877 => (x"00",x"00",x"2e",x"d2"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"13",x"43"),
  1880 => (x"00",x"00",x"2e",x"f0"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"16",x"5d"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"00",x"00",x"13",x"f7"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"db",x"86",x"fc",x"1e"),
  1889 => (x"fc",x"7e",x"70",x"87"),
  1890 => (x"1e",x"4f",x"26",x"8e"),
  1891 => (x"c0",x"48",x"f0",x"fe"),
  1892 => (x"79",x"09",x"cd",x"78"),
  1893 => (x"1e",x"4f",x"26",x"09"),
  1894 => (x"49",x"c0",x"f6",x"c1"),
  1895 => (x"4f",x"26",x"87",x"ed"),
  1896 => (x"bf",x"f0",x"fe",x"1e"),
  1897 => (x"1e",x"4f",x"26",x"48"),
  1898 => (x"c1",x"48",x"f0",x"fe"),
  1899 => (x"1e",x"4f",x"26",x"78"),
  1900 => (x"c0",x"48",x"f0",x"fe"),
  1901 => (x"1e",x"4f",x"26",x"78"),
  1902 => (x"52",x"c0",x"4a",x"71"),
  1903 => (x"0e",x"4f",x"26",x"51"),
  1904 => (x"5d",x"5c",x"5b",x"5e"),
  1905 => (x"71",x"86",x"f4",x"0e"),
  1906 => (x"7e",x"6d",x"97",x"4d"),
  1907 => (x"97",x"4c",x"a5",x"c1"),
  1908 => (x"a6",x"c8",x"48",x"6c"),
  1909 => (x"c4",x"48",x"6e",x"58"),
  1910 => (x"c5",x"05",x"a8",x"66"),
  1911 => (x"c0",x"48",x"ff",x"87"),
  1912 => (x"ca",x"ff",x"87",x"e6"),
  1913 => (x"49",x"a5",x"c2",x"87"),
  1914 => (x"71",x"4b",x"6c",x"97"),
  1915 => (x"6b",x"97",x"4b",x"a3"),
  1916 => (x"7e",x"6c",x"97",x"4b"),
  1917 => (x"80",x"c1",x"48",x"6e"),
  1918 => (x"c7",x"58",x"a6",x"c8"),
  1919 => (x"58",x"a6",x"cc",x"98"),
  1920 => (x"fe",x"7c",x"97",x"70"),
  1921 => (x"48",x"73",x"87",x"e1"),
  1922 => (x"4d",x"26",x"8e",x"f4"),
  1923 => (x"4b",x"26",x"4c",x"26"),
  1924 => (x"5e",x"0e",x"4f",x"26"),
  1925 => (x"f4",x"0e",x"5c",x"5b"),
  1926 => (x"d8",x"4c",x"71",x"86"),
  1927 => (x"ff",x"c3",x"4a",x"66"),
  1928 => (x"4b",x"a4",x"c2",x"9a"),
  1929 => (x"73",x"49",x"6c",x"97"),
  1930 => (x"51",x"72",x"49",x"a1"),
  1931 => (x"6e",x"7e",x"6c",x"97"),
  1932 => (x"c8",x"80",x"c1",x"48"),
  1933 => (x"98",x"c7",x"58",x"a6"),
  1934 => (x"70",x"58",x"a6",x"cc"),
  1935 => (x"26",x"8e",x"f4",x"54"),
  1936 => (x"26",x"4b",x"26",x"4c"),
  1937 => (x"86",x"fc",x"1e",x"4f"),
  1938 => (x"e0",x"87",x"e4",x"fd"),
  1939 => (x"c0",x"49",x"4a",x"bf"),
  1940 => (x"02",x"99",x"c0",x"e0"),
  1941 => (x"1e",x"72",x"87",x"cb"),
  1942 => (x"49",x"d0",x"fc",x"c2"),
  1943 => (x"c4",x"87",x"f3",x"fe"),
  1944 => (x"87",x"fc",x"fc",x"86"),
  1945 => (x"fe",x"fc",x"7e",x"70"),
  1946 => (x"26",x"8e",x"fc",x"87"),
  1947 => (x"fc",x"c2",x"1e",x"4f"),
  1948 => (x"c2",x"fd",x"49",x"d0"),
  1949 => (x"c5",x"f9",x"c1",x"87"),
  1950 => (x"87",x"cf",x"fc",x"49"),
  1951 => (x"26",x"87",x"ed",x"c3"),
  1952 => (x"5b",x"5e",x"0e",x"4f"),
  1953 => (x"fc",x"0e",x"5d",x"5c"),
  1954 => (x"ff",x"7e",x"71",x"86"),
  1955 => (x"fc",x"c2",x"4d",x"d4"),
  1956 => (x"ea",x"fc",x"49",x"d0"),
  1957 => (x"c0",x"4b",x"70",x"87"),
  1958 => (x"c2",x"04",x"ab",x"b7"),
  1959 => (x"f0",x"c3",x"87",x"f8"),
  1960 => (x"87",x"c9",x"05",x"ab"),
  1961 => (x"48",x"e4",x"fd",x"c1"),
  1962 => (x"d9",x"c2",x"78",x"c1"),
  1963 => (x"ab",x"e0",x"c3",x"87"),
  1964 => (x"c1",x"87",x"c9",x"05"),
  1965 => (x"c1",x"48",x"e8",x"fd"),
  1966 => (x"87",x"ca",x"c2",x"78"),
  1967 => (x"bf",x"e8",x"fd",x"c1"),
  1968 => (x"c2",x"87",x"c6",x"02"),
  1969 => (x"c2",x"4c",x"a3",x"c0"),
  1970 => (x"c1",x"4c",x"73",x"87"),
  1971 => (x"02",x"bf",x"e4",x"fd"),
  1972 => (x"74",x"87",x"e0",x"c0"),
  1973 => (x"29",x"b7",x"c4",x"49"),
  1974 => (x"c0",x"ff",x"c1",x"91"),
  1975 => (x"cf",x"4a",x"74",x"81"),
  1976 => (x"c1",x"92",x"c2",x"9a"),
  1977 => (x"70",x"30",x"72",x"48"),
  1978 => (x"72",x"ba",x"ff",x"4a"),
  1979 => (x"70",x"98",x"69",x"48"),
  1980 => (x"74",x"87",x"db",x"79"),
  1981 => (x"29",x"b7",x"c4",x"49"),
  1982 => (x"c0",x"ff",x"c1",x"91"),
  1983 => (x"cf",x"4a",x"74",x"81"),
  1984 => (x"c3",x"92",x"c2",x"9a"),
  1985 => (x"70",x"30",x"72",x"48"),
  1986 => (x"b0",x"69",x"48",x"4a"),
  1987 => (x"05",x"6e",x"79",x"70"),
  1988 => (x"ff",x"87",x"e7",x"c0"),
  1989 => (x"e1",x"c8",x"48",x"d0"),
  1990 => (x"c1",x"7d",x"c5",x"78"),
  1991 => (x"02",x"bf",x"e8",x"fd"),
  1992 => (x"e0",x"c3",x"87",x"c3"),
  1993 => (x"e4",x"fd",x"c1",x"7d"),
  1994 => (x"87",x"c3",x"02",x"bf"),
  1995 => (x"73",x"7d",x"f0",x"c3"),
  1996 => (x"48",x"d0",x"ff",x"7d"),
  1997 => (x"c0",x"78",x"e1",x"c8"),
  1998 => (x"fd",x"c1",x"78",x"e0"),
  1999 => (x"78",x"c0",x"48",x"e8"),
  2000 => (x"48",x"e4",x"fd",x"c1"),
  2001 => (x"fc",x"c2",x"78",x"c0"),
  2002 => (x"f2",x"f9",x"49",x"d0"),
  2003 => (x"c0",x"4b",x"70",x"87"),
  2004 => (x"fd",x"03",x"ab",x"b7"),
  2005 => (x"48",x"c0",x"87",x"c8"),
  2006 => (x"4d",x"26",x"8e",x"fc"),
  2007 => (x"4b",x"26",x"4c",x"26"),
  2008 => (x"00",x"00",x"4f",x"26"),
  2009 => (x"00",x"00",x"00",x"00"),
  2010 => (x"00",x"00",x"00",x"00"),
  2011 => (x"72",x"4a",x"c0",x"1e"),
  2012 => (x"c1",x"91",x"c4",x"49"),
  2013 => (x"c0",x"81",x"c0",x"ff"),
  2014 => (x"d0",x"82",x"c1",x"79"),
  2015 => (x"ee",x"04",x"aa",x"b7"),
  2016 => (x"0e",x"4f",x"26",x"87"),
  2017 => (x"5d",x"5c",x"5b",x"5e"),
  2018 => (x"f8",x"4d",x"71",x"0e"),
  2019 => (x"4a",x"75",x"87",x"e1"),
  2020 => (x"92",x"2a",x"b7",x"c4"),
  2021 => (x"82",x"c0",x"ff",x"c1"),
  2022 => (x"9c",x"cf",x"4c",x"75"),
  2023 => (x"49",x"6a",x"94",x"c2"),
  2024 => (x"c3",x"2b",x"74",x"4b"),
  2025 => (x"74",x"48",x"c2",x"9b"),
  2026 => (x"ff",x"4c",x"70",x"30"),
  2027 => (x"71",x"48",x"74",x"bc"),
  2028 => (x"f7",x"7a",x"70",x"98"),
  2029 => (x"48",x"73",x"87",x"f1"),
  2030 => (x"4c",x"26",x"4d",x"26"),
  2031 => (x"4f",x"26",x"4b",x"26"),
  2032 => (x"00",x"00",x"00",x"00"),
  2033 => (x"00",x"00",x"00",x"00"),
  2034 => (x"00",x"00",x"00",x"00"),
  2035 => (x"00",x"00",x"00",x"00"),
  2036 => (x"00",x"00",x"00",x"00"),
  2037 => (x"00",x"00",x"00",x"00"),
  2038 => (x"00",x"00",x"00",x"00"),
  2039 => (x"00",x"00",x"00",x"00"),
  2040 => (x"00",x"00",x"00",x"00"),
  2041 => (x"00",x"00",x"00",x"00"),
  2042 => (x"00",x"00",x"00",x"00"),
  2043 => (x"00",x"00",x"00",x"00"),
  2044 => (x"00",x"00",x"00",x"00"),
  2045 => (x"00",x"00",x"00",x"00"),
  2046 => (x"00",x"00",x"00",x"00"),
  2047 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

